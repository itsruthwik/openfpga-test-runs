//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug 20 23:29:10 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__5_ -----
module sb_1__5_(pReset,
                prog_clk,
                chany_top_in,
                chanx_right_in,
                chany_bottom_in,
                chanx_left_in,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:104] chany_top_in;
//----- INPUT PORTS -----
input [0:104] chanx_right_in;
//----- INPUT PORTS -----
input [0:104] chany_bottom_in;
//----- INPUT PORTS -----
input [0:104] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:104] chany_top_out;
//----- OUTPUT PORTS -----
output [0:104] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:104] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:104] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:5] mux_2level_tapbuf_size6_0_sram;
wire [0:5] mux_2level_tapbuf_size6_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_1_sram;
wire [0:5] mux_2level_tapbuf_size6_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_1_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_10_sram;
wire [0:5] mux_2level_tapbuf_size7_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_11_sram;
wire [0:5] mux_2level_tapbuf_size7_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_12_sram;
wire [0:5] mux_2level_tapbuf_size7_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_13_sram;
wire [0:5] mux_2level_tapbuf_size7_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_14_sram;
wire [0:5] mux_2level_tapbuf_size7_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_15_sram;
wire [0:5] mux_2level_tapbuf_size7_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_16_sram;
wire [0:5] mux_2level_tapbuf_size7_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_17_sram;
wire [0:5] mux_2level_tapbuf_size7_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_18_sram;
wire [0:5] mux_2level_tapbuf_size7_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_19_sram;
wire [0:5] mux_2level_tapbuf_size7_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_4_sram;
wire [0:5] mux_2level_tapbuf_size7_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_5_sram;
wire [0:5] mux_2level_tapbuf_size7_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_6_sram;
wire [0:5] mux_2level_tapbuf_size7_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_7_sram;
wire [0:5] mux_2level_tapbuf_size7_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_8_sram;
wire [0:5] mux_2level_tapbuf_size7_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_9_sram;
wire [0:5] mux_2level_tapbuf_size7_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_16_sram;
wire [0:5] mux_2level_tapbuf_size8_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_17_sram;
wire [0:5] mux_2level_tapbuf_size8_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_18_sram;
wire [0:5] mux_2level_tapbuf_size8_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_19_sram;
wire [0:5] mux_2level_tapbuf_size8_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_20_sram;
wire [0:5] mux_2level_tapbuf_size8_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_21_sram;
wire [0:5] mux_2level_tapbuf_size8_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_22_sram;
wire [0:5] mux_2level_tapbuf_size8_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_23_sram;
wire [0:5] mux_2level_tapbuf_size8_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_24_sram;
wire [0:5] mux_2level_tapbuf_size8_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_25_sram;
wire [0:5] mux_2level_tapbuf_size8_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_26_sram;
wire [0:5] mux_2level_tapbuf_size8_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_27_sram;
wire [0:5] mux_2level_tapbuf_size8_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_28_sram;
wire [0:5] mux_2level_tapbuf_size8_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_29_sram;
wire [0:5] mux_2level_tapbuf_size8_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_30_sram;
wire [0:5] mux_2level_tapbuf_size8_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_31_sram;
wire [0:5] mux_2level_tapbuf_size8_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_32_sram;
wire [0:5] mux_2level_tapbuf_size8_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_33_sram;
wire [0:5] mux_2level_tapbuf_size8_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_34_sram;
wire [0:5] mux_2level_tapbuf_size8_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_35_sram;
wire [0:5] mux_2level_tapbuf_size8_35_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_36_sram;
wire [0:5] mux_2level_tapbuf_size8_36_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_37_sram;
wire [0:5] mux_2level_tapbuf_size8_37_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_38_sram;
wire [0:5] mux_2level_tapbuf_size8_38_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_39_sram;
wire [0:5] mux_2level_tapbuf_size8_39_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_40_sram;
wire [0:5] mux_2level_tapbuf_size8_40_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_41_sram;
wire [0:5] mux_2level_tapbuf_size8_41_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_42_sram;
wire [0:5] mux_2level_tapbuf_size8_42_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_43_sram;
wire [0:5] mux_2level_tapbuf_size8_43_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_44_sram;
wire [0:5] mux_2level_tapbuf_size8_44_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_45_sram;
wire [0:5] mux_2level_tapbuf_size8_45_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_46_sram;
wire [0:5] mux_2level_tapbuf_size8_46_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_47_sram;
wire [0:5] mux_2level_tapbuf_size8_47_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_48_sram;
wire [0:5] mux_2level_tapbuf_size8_48_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_49_sram;
wire [0:5] mux_2level_tapbuf_size8_49_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_50_sram;
wire [0:5] mux_2level_tapbuf_size8_50_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_51_sram;
wire [0:5] mux_2level_tapbuf_size8_51_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_52_sram;
wire [0:5] mux_2level_tapbuf_size8_52_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_53_sram;
wire [0:5] mux_2level_tapbuf_size8_53_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_54_sram;
wire [0:5] mux_2level_tapbuf_size8_54_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_55_sram;
wire [0:5] mux_2level_tapbuf_size8_55_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_56_sram;
wire [0:5] mux_2level_tapbuf_size8_56_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_57_sram;
wire [0:5] mux_2level_tapbuf_size8_57_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_58_sram;
wire [0:5] mux_2level_tapbuf_size8_58_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_59_sram;
wire [0:5] mux_2level_tapbuf_size8_59_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_60_sram;
wire [0:5] mux_2level_tapbuf_size8_60_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_61_sram;
wire [0:5] mux_2level_tapbuf_size8_61_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_62_sram;
wire [0:5] mux_2level_tapbuf_size8_62_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_63_sram;
wire [0:5] mux_2level_tapbuf_size8_63_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_64_sram;
wire [0:5] mux_2level_tapbuf_size8_64_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_65_sram;
wire [0:5] mux_2level_tapbuf_size8_65_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_66_sram;
wire [0:5] mux_2level_tapbuf_size8_66_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_67_sram;
wire [0:5] mux_2level_tapbuf_size8_67_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_68_sram;
wire [0:5] mux_2level_tapbuf_size8_68_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_69_sram;
wire [0:5] mux_2level_tapbuf_size8_69_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_70_sram;
wire [0:5] mux_2level_tapbuf_size8_70_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_71_sram;
wire [0:5] mux_2level_tapbuf_size8_71_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_72_sram;
wire [0:5] mux_2level_tapbuf_size8_72_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_73_sram;
wire [0:5] mux_2level_tapbuf_size8_73_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_74_sram;
wire [0:5] mux_2level_tapbuf_size8_74_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_75_sram;
wire [0:5] mux_2level_tapbuf_size8_75_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_76_sram;
wire [0:5] mux_2level_tapbuf_size8_76_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_77_sram;
wire [0:5] mux_2level_tapbuf_size8_77_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_78_sram;
wire [0:5] mux_2level_tapbuf_size8_78_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_79_sram;
wire [0:5] mux_2level_tapbuf_size8_79_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_80_sram;
wire [0:5] mux_2level_tapbuf_size8_80_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_81_sram;
wire [0:5] mux_2level_tapbuf_size8_81_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_82_sram;
wire [0:5] mux_2level_tapbuf_size8_82_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_83_sram;
wire [0:5] mux_2level_tapbuf_size8_83_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_84_sram;
wire [0:5] mux_2level_tapbuf_size8_84_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_85_sram;
wire [0:5] mux_2level_tapbuf_size8_85_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size8 mux_top_track_0 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[37], chanx_right_in[73], chanx_left_in[0], chanx_left_in[3], chanx_left_in[36], chanx_left_in[72]}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size8 mux_top_track_32 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[42], chanx_right_in[78], chanx_left_in[30], chanx_left_in[66], chanx_left_in[95], chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size8 mux_top_track_40 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[44], chanx_right_in[80], chanx_left_in[29], chanx_left_in[65], chanx_left_in[91], chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size8 mux_top_track_48 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[45], chanx_right_in[81], chanx_left_in[28], chanx_left_in[64], chanx_left_in[87], chanx_left_in[100]}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size8 mux_top_track_56 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[46], chanx_right_in[82], chanx_left_in[26], chanx_left_in[62], chanx_left_in[83], chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size8 mux_top_track_64 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[48], chanx_right_in[84], chanx_left_in[25], chanx_left_in[61], chanx_left_in[79], chanx_left_in[97]}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size8 mux_top_track_72 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[49], chanx_right_in[85], chanx_left_in[24], chanx_left_in[60], chanx_left_in[75], chanx_left_in[96]}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size8 mux_top_track_80 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[50], chanx_right_in[86], chanx_left_in[22], chanx_left_in[58], chanx_left_in[71], chanx_left_in[94]}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size8 mux_top_track_88 (
		.in({chanx_right_in[16], chanx_right_in[51:52], chanx_right_in[88], chanx_left_in[21], chanx_left_in[57], chanx_left_in[67], chanx_left_in[93]}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size8 mux_top_track_96 (
		.in({chanx_right_in[17], chanx_right_in[53], chanx_right_in[55], chanx_right_in[89], chanx_left_in[20], chanx_left_in[56], chanx_left_in[63], chanx_left_in[92]}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size8 mux_top_track_104 (
		.in({chanx_right_in[18], chanx_right_in[54], chanx_right_in[59], chanx_right_in[90], chanx_left_in[18], chanx_left_in[54], chanx_left_in[59], chanx_left_in[90]}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size8 mux_top_track_112 (
		.in({chanx_right_in[20], chanx_right_in[56], chanx_right_in[63], chanx_right_in[92], chanx_left_in[17], chanx_left_in[53], chanx_left_in[55], chanx_left_in[89]}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size8 mux_top_track_120 (
		.in({chanx_right_in[21], chanx_right_in[57], chanx_right_in[67], chanx_right_in[93], chanx_left_in[16], chanx_left_in[51:52], chanx_left_in[88]}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size8 mux_top_track_128 (
		.in({chanx_right_in[22], chanx_right_in[58], chanx_right_in[71], chanx_right_in[94], chanx_left_in[14], chanx_left_in[47], chanx_left_in[50], chanx_left_in[86]}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size8 mux_top_track_136 (
		.in({chanx_right_in[24], chanx_right_in[60], chanx_right_in[75], chanx_right_in[96], chanx_left_in[13], chanx_left_in[43], chanx_left_in[49], chanx_left_in[85]}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size8 mux_top_track_144 (
		.in({chanx_right_in[25], chanx_right_in[61], chanx_right_in[79], chanx_right_in[97], chanx_left_in[12], chanx_left_in[39], chanx_left_in[48], chanx_left_in[84]}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size8 mux_top_track_152 (
		.in({chanx_right_in[26], chanx_right_in[62], chanx_right_in[83], chanx_right_in[98], chanx_left_in[10], chanx_left_in[35], chanx_left_in[46], chanx_left_in[82]}),
		.sram(mux_2level_tapbuf_size8_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_16_sram_inv[0:5]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size8 mux_top_track_160 (
		.in({chanx_right_in[28], chanx_right_in[64], chanx_right_in[87], chanx_right_in[100], chanx_left_in[9], chanx_left_in[31], chanx_left_in[45], chanx_left_in[81]}),
		.sram(mux_2level_tapbuf_size8_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_17_sram_inv[0:5]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size8 mux_top_track_168 (
		.in({chanx_right_in[29], chanx_right_in[65], chanx_right_in[91], chanx_right_in[101], chanx_left_in[8], chanx_left_in[27], chanx_left_in[44], chanx_left_in[80]}),
		.sram(mux_2level_tapbuf_size8_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_18_sram_inv[0:5]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size8 mux_top_track_176 (
		.in({chanx_right_in[30], chanx_right_in[66], chanx_right_in[95], chanx_right_in[102], chanx_left_in[6], chanx_left_in[23], chanx_left_in[42], chanx_left_in[78]}),
		.sram(mux_2level_tapbuf_size8_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_19_sram_inv[0:5]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size8 mux_top_track_208 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[36], chanx_right_in[72], chanx_left_in[1], chanx_left_in[7], chanx_left_in[37], chanx_left_in[73]}),
		.sram(mux_2level_tapbuf_size8_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_20_sram_inv[0:5]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size8 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[37], chany_top_in[73], chany_bottom_in[30], chany_bottom_in[66], chany_bottom_in[95], chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size8_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_21_sram_inv[0:5]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size8 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[38], chany_top_in[74], chany_bottom_in[29], chany_bottom_in[65], chany_bottom_in[91], chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size8_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_22_sram_inv[0:5]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size8 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[40], chany_top_in[76], chany_bottom_in[28], chany_bottom_in[64], chany_bottom_in[87], chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size8_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_23_sram_inv[0:5]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size8 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[41], chany_top_in[77], chany_bottom_in[26], chany_bottom_in[62], chany_bottom_in[83], chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size8_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_24_sram_inv[0:5]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size8 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[42], chany_top_in[78], chany_bottom_in[25], chany_bottom_in[61], chany_bottom_in[79], chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size8_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_25_sram_inv[0:5]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size8 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[44], chany_top_in[80], chany_bottom_in[24], chany_bottom_in[60], chany_bottom_in[75], chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size8_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_26_sram_inv[0:5]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size8 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[45], chany_top_in[81], chany_bottom_in[22], chany_bottom_in[58], chany_bottom_in[71], chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size8_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_27_sram_inv[0:5]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size8 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[46], chany_top_in[82], chany_bottom_in[21], chany_bottom_in[57], chany_bottom_in[67], chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size8_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_28_sram_inv[0:5]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size8 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[48], chany_top_in[84], chany_bottom_in[20], chany_bottom_in[56], chany_bottom_in[63], chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size8_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_29_sram_inv[0:5]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size8 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[49], chany_top_in[85], chany_bottom_in[18], chany_bottom_in[54], chany_bottom_in[59], chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size8_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_30_sram_inv[0:5]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size8 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[50], chany_top_in[86], chany_bottom_in[17], chany_bottom_in[53], chany_bottom_in[55], chany_bottom_in[89]}),
		.sram(mux_2level_tapbuf_size8_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_31_sram_inv[0:5]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size8 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51:52], chany_top_in[88], chany_bottom_in[16], chany_bottom_in[51:52], chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size8_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_32_sram_inv[0:5]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size8 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[53], chany_top_in[55], chany_top_in[89], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[50], chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size8_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_33_sram_inv[0:5]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size8 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[54], chany_top_in[59], chany_top_in[90], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[49], chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size8_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_34_sram_inv[0:5]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size8 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[56], chany_top_in[63], chany_top_in[92], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[48], chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size8_35_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_35_sram_inv[0:5]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size8 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[57], chany_top_in[67], chany_top_in[93], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[46], chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size8_36_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_36_sram_inv[0:5]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size8 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[58], chany_top_in[71], chany_top_in[94], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[45], chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size8_37_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_37_sram_inv[0:5]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size8 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[60], chany_top_in[75], chany_top_in[96], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[44], chany_bottom_in[80]}),
		.sram(mux_2level_tapbuf_size8_38_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_38_sram_inv[0:5]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size8 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[61], chany_top_in[79], chany_top_in[97], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[42], chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size8_39_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_39_sram_inv[0:5]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size8 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[62], chany_top_in[83], chany_top_in[98], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[41], chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size8_40_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_40_sram_inv[0:5]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size8 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[64], chany_top_in[87], chany_top_in[100], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[40], chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size8_41_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_41_sram_inv[0:5]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size8 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[65], chany_top_in[91], chany_top_in[101], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[38], chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size8_42_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_42_sram_inv[0:5]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size8 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[66], chany_top_in[95], chany_top_in[102], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size8_43_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_43_sram_inv[0:5]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size8 mux_bottom_track_17 (
		.in({chanx_right_in[30], chanx_right_in[66], chanx_right_in[95], chanx_right_in[102], chanx_left_in[4], chanx_left_in[15], chanx_left_in[40], chanx_left_in[76]}),
		.sram(mux_2level_tapbuf_size8_44_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_44_sram_inv[0:5]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size8 mux_bottom_track_25 (
		.in({chanx_right_in[29], chanx_right_in[65], chanx_right_in[91], chanx_right_in[101], chanx_left_in[5], chanx_left_in[19], chanx_left_in[41], chanx_left_in[77]}),
		.sram(mux_2level_tapbuf_size8_45_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_45_sram_inv[0:5]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size8 mux_bottom_track_33 (
		.in({chanx_right_in[28], chanx_right_in[64], chanx_right_in[87], chanx_right_in[100], chanx_left_in[6], chanx_left_in[23], chanx_left_in[42], chanx_left_in[78]}),
		.sram(mux_2level_tapbuf_size8_46_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_46_sram_inv[0:5]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size8 mux_bottom_track_41 (
		.in({chanx_right_in[26], chanx_right_in[62], chanx_right_in[83], chanx_right_in[98], chanx_left_in[8], chanx_left_in[27], chanx_left_in[44], chanx_left_in[80]}),
		.sram(mux_2level_tapbuf_size8_47_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_47_sram_inv[0:5]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size8 mux_bottom_track_49 (
		.in({chanx_right_in[25], chanx_right_in[61], chanx_right_in[79], chanx_right_in[97], chanx_left_in[9], chanx_left_in[31], chanx_left_in[45], chanx_left_in[81]}),
		.sram(mux_2level_tapbuf_size8_48_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_48_sram_inv[0:5]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size8 mux_bottom_track_57 (
		.in({chanx_right_in[24], chanx_right_in[60], chanx_right_in[75], chanx_right_in[96], chanx_left_in[10], chanx_left_in[35], chanx_left_in[46], chanx_left_in[82]}),
		.sram(mux_2level_tapbuf_size8_49_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_49_sram_inv[0:5]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size8 mux_bottom_track_65 (
		.in({chanx_right_in[22], chanx_right_in[58], chanx_right_in[71], chanx_right_in[94], chanx_left_in[12], chanx_left_in[39], chanx_left_in[48], chanx_left_in[84]}),
		.sram(mux_2level_tapbuf_size8_50_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_50_sram_inv[0:5]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size8 mux_bottom_track_73 (
		.in({chanx_right_in[21], chanx_right_in[57], chanx_right_in[67], chanx_right_in[93], chanx_left_in[13], chanx_left_in[43], chanx_left_in[49], chanx_left_in[85]}),
		.sram(mux_2level_tapbuf_size8_51_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_51_sram_inv[0:5]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size8 mux_bottom_track_81 (
		.in({chanx_right_in[20], chanx_right_in[56], chanx_right_in[63], chanx_right_in[92], chanx_left_in[14], chanx_left_in[47], chanx_left_in[50], chanx_left_in[86]}),
		.sram(mux_2level_tapbuf_size8_52_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_52_sram_inv[0:5]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size8 mux_bottom_track_89 (
		.in({chanx_right_in[18], chanx_right_in[54], chanx_right_in[59], chanx_right_in[90], chanx_left_in[16], chanx_left_in[51:52], chanx_left_in[88]}),
		.sram(mux_2level_tapbuf_size8_53_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_53_sram_inv[0:5]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size8 mux_bottom_track_97 (
		.in({chanx_right_in[17], chanx_right_in[53], chanx_right_in[55], chanx_right_in[89], chanx_left_in[17], chanx_left_in[53], chanx_left_in[55], chanx_left_in[89]}),
		.sram(mux_2level_tapbuf_size8_54_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_54_sram_inv[0:5]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size8 mux_bottom_track_105 (
		.in({chanx_right_in[16], chanx_right_in[51:52], chanx_right_in[88], chanx_left_in[18], chanx_left_in[54], chanx_left_in[59], chanx_left_in[90]}),
		.sram(mux_2level_tapbuf_size8_55_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_55_sram_inv[0:5]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size8 mux_bottom_track_113 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[50], chanx_right_in[86], chanx_left_in[20], chanx_left_in[56], chanx_left_in[63], chanx_left_in[92]}),
		.sram(mux_2level_tapbuf_size8_56_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_56_sram_inv[0:5]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size8 mux_bottom_track_121 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[49], chanx_right_in[85], chanx_left_in[21], chanx_left_in[57], chanx_left_in[67], chanx_left_in[93]}),
		.sram(mux_2level_tapbuf_size8_57_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_57_sram_inv[0:5]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size8 mux_bottom_track_129 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[48], chanx_right_in[84], chanx_left_in[22], chanx_left_in[58], chanx_left_in[71], chanx_left_in[94]}),
		.sram(mux_2level_tapbuf_size8_58_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_58_sram_inv[0:5]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size8 mux_bottom_track_137 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[46], chanx_right_in[82], chanx_left_in[24], chanx_left_in[60], chanx_left_in[75], chanx_left_in[96]}),
		.sram(mux_2level_tapbuf_size8_59_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_59_sram_inv[0:5]),
		.out(chany_bottom_out[68]));

	mux_2level_tapbuf_size8 mux_bottom_track_145 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[45], chanx_right_in[81], chanx_left_in[25], chanx_left_in[61], chanx_left_in[79], chanx_left_in[97]}),
		.sram(mux_2level_tapbuf_size8_60_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_60_sram_inv[0:5]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size8 mux_bottom_track_153 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[44], chanx_right_in[80], chanx_left_in[26], chanx_left_in[62], chanx_left_in[83], chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size8_61_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_61_sram_inv[0:5]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size8 mux_bottom_track_161 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[42], chanx_right_in[78], chanx_left_in[28], chanx_left_in[64], chanx_left_in[87], chanx_left_in[100]}),
		.sram(mux_2level_tapbuf_size8_62_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_62_sram_inv[0:5]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size8 mux_bottom_track_169 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[41], chanx_right_in[77], chanx_left_in[29], chanx_left_in[65], chanx_left_in[91], chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size8_63_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_63_sram_inv[0:5]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size8 mux_bottom_track_177 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[40], chanx_right_in[76], chanx_left_in[30], chanx_left_in[66], chanx_left_in[95], chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size8_64_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_64_sram_inv[0:5]),
		.out(chany_bottom_out[88]));

	mux_2level_tapbuf_size8 mux_left_track_33 (
		.in({chany_top_in[30], chany_top_in[66], chany_top_in[95], chany_top_in[102], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[40], chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size8_65_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_65_sram_inv[0:5]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size8 mux_left_track_41 (
		.in({chany_top_in[29], chany_top_in[65], chany_top_in[91], chany_top_in[101], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[41], chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size8_66_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_66_sram_inv[0:5]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size8 mux_left_track_49 (
		.in({chany_top_in[28], chany_top_in[64], chany_top_in[87], chany_top_in[100], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[42], chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size8_67_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_67_sram_inv[0:5]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size8 mux_left_track_57 (
		.in({chany_top_in[26], chany_top_in[62], chany_top_in[83], chany_top_in[98], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[44], chany_bottom_in[80]}),
		.sram(mux_2level_tapbuf_size8_68_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_68_sram_inv[0:5]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size8 mux_left_track_65 (
		.in({chany_top_in[25], chany_top_in[61], chany_top_in[79], chany_top_in[97], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[45], chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size8_69_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_69_sram_inv[0:5]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size8 mux_left_track_73 (
		.in({chany_top_in[24], chany_top_in[60], chany_top_in[75], chany_top_in[96], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[46], chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size8_70_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_70_sram_inv[0:5]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size8 mux_left_track_81 (
		.in({chany_top_in[22], chany_top_in[58], chany_top_in[71], chany_top_in[94], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[48], chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size8_71_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_71_sram_inv[0:5]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size8 mux_left_track_89 (
		.in({chany_top_in[21], chany_top_in[57], chany_top_in[67], chany_top_in[93], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[49], chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size8_72_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_72_sram_inv[0:5]),
		.out(chanx_left_out[44]));

	mux_2level_tapbuf_size8 mux_left_track_97 (
		.in({chany_top_in[20], chany_top_in[56], chany_top_in[63], chany_top_in[92], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[50], chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size8_73_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_73_sram_inv[0:5]),
		.out(chanx_left_out[48]));

	mux_2level_tapbuf_size8 mux_left_track_105 (
		.in({chany_top_in[18], chany_top_in[54], chany_top_in[59], chany_top_in[90], chany_bottom_in[16], chany_bottom_in[51:52], chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size8_74_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_74_sram_inv[0:5]),
		.out(chanx_left_out[52]));

	mux_2level_tapbuf_size8 mux_left_track_113 (
		.in({chany_top_in[17], chany_top_in[53], chany_top_in[55], chany_top_in[89], chany_bottom_in[17], chany_bottom_in[53], chany_bottom_in[55], chany_bottom_in[89]}),
		.sram(mux_2level_tapbuf_size8_75_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_75_sram_inv[0:5]),
		.out(chanx_left_out[56]));

	mux_2level_tapbuf_size8 mux_left_track_121 (
		.in({chany_top_in[16], chany_top_in[51:52], chany_top_in[88], chany_bottom_in[18], chany_bottom_in[54], chany_bottom_in[59], chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size8_76_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_76_sram_inv[0:5]),
		.out(chanx_left_out[60]));

	mux_2level_tapbuf_size8 mux_left_track_129 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[50], chany_top_in[86], chany_bottom_in[20], chany_bottom_in[56], chany_bottom_in[63], chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size8_77_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_77_sram_inv[0:5]),
		.out(chanx_left_out[64]));

	mux_2level_tapbuf_size8 mux_left_track_137 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[49], chany_top_in[85], chany_bottom_in[21], chany_bottom_in[57], chany_bottom_in[67], chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size8_78_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_78_sram_inv[0:5]),
		.out(chanx_left_out[68]));

	mux_2level_tapbuf_size8 mux_left_track_145 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[48], chany_top_in[84], chany_bottom_in[22], chany_bottom_in[58], chany_bottom_in[71], chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size8_79_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_79_sram_inv[0:5]),
		.out(chanx_left_out[72]));

	mux_2level_tapbuf_size8 mux_left_track_153 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[46], chany_top_in[82], chany_bottom_in[24], chany_bottom_in[60], chany_bottom_in[75], chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size8_80_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_80_sram_inv[0:5]),
		.out(chanx_left_out[76]));

	mux_2level_tapbuf_size8 mux_left_track_161 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[45], chany_top_in[81], chany_bottom_in[25], chany_bottom_in[61], chany_bottom_in[79], chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size8_81_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_81_sram_inv[0:5]),
		.out(chanx_left_out[80]));

	mux_2level_tapbuf_size8 mux_left_track_169 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[44], chany_top_in[80], chany_bottom_in[26], chany_bottom_in[62], chany_bottom_in[83], chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size8_82_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_82_sram_inv[0:5]),
		.out(chanx_left_out[84]));

	mux_2level_tapbuf_size8 mux_left_track_177 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[42], chany_top_in[78], chany_bottom_in[28], chany_bottom_in[64], chany_bottom_in[87], chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size8_83_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_83_sram_inv[0:5]),
		.out(chanx_left_out[88]));

	mux_2level_tapbuf_size8 mux_left_track_185 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[41], chany_top_in[77], chany_bottom_in[29], chany_bottom_in[65], chany_bottom_in[91], chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size8_84_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_84_sram_inv[0:5]),
		.out(chanx_left_out[92]));

	mux_2level_tapbuf_size8 mux_left_track_193 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[40], chany_top_in[76], chany_bottom_in[30], chany_bottom_in[66], chany_bottom_in[95], chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size8_85_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_85_sram_inv[0:5]),
		.out(chanx_left_out[96]));

	mux_2level_tapbuf_size8_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_16_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_17_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_18_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_19_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_20_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_21_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_22_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_23_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_24_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_25_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_26_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_27_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_28_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_29_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_30_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_31_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_32_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_33_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_34_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_35_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_35_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_36_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_36_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_37_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_37_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_38_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_38_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_39_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_39_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_40_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_40_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_41_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_41_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_42_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_42_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_43_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_43_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_44_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_44_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_45_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_45_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_46_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_46_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_47_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_47_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_48_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_48_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_49_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_49_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_50_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_50_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_51_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_51_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_52_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_52_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_53_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_53_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_54_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_54_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_55_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_55_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_56_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_56_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_57_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_57_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_58_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_58_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_59_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_59_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_60_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_60_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_61_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_61_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_62_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_62_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_63_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_63_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_64_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_64_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_65_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_65_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_66_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_66_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_67_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_67_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_68_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_68_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_69_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_69_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_70_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_70_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_71_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_71_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_72_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_72_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_73_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_73_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_74_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_74_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_75_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_75_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_76_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_76_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_77_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_77_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_78_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_78_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_79_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_79_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_80_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_80_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_81_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_81_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_82_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_82_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_83_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_83_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_84_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_84_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_85_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_85_sram_inv[0:5]));

	mux_2level_tapbuf_size7 mux_top_track_8 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[38], chanx_right_in[74], chanx_left_in[34], chanx_left_in[70], chanx_left_in[104]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size7 mux_top_track_16 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[40], chanx_right_in[76], chanx_left_in[33], chanx_left_in[69], chanx_left_in[103]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size7 mux_top_track_24 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[41], chanx_right_in[77], chanx_left_in[32], chanx_left_in[68], chanx_left_in[99]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size7 mux_top_track_184 (
		.in({chanx_right_in[32], chanx_right_in[68], chanx_right_in[99], chanx_left_in[5], chanx_left_in[19], chanx_left_in[41], chanx_left_in[77]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size7 mux_top_track_192 (
		.in({chanx_right_in[33], chanx_right_in[69], chanx_right_in[103], chanx_left_in[4], chanx_left_in[15], chanx_left_in[40], chanx_left_in[76]}),
		.sram(mux_2level_tapbuf_size7_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_4_sram_inv[0:5]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size7 mux_top_track_200 (
		.in({chanx_right_in[34], chanx_right_in[70], chanx_right_in[104], chanx_left_in[2], chanx_left_in[11], chanx_left_in[38], chanx_left_in[74]}),
		.sram(mux_2level_tapbuf_size7_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_5_sram_inv[0:5]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size7 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[36], chany_top_in[72], chany_bottom_in[32], chany_bottom_in[68], chany_bottom_in[99]}),
		.sram(mux_2level_tapbuf_size7_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_6_sram_inv[0:5]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size7 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[68], chany_top_in[99], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[36], chany_bottom_in[72]}),
		.sram(mux_2level_tapbuf_size7_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_7_sram_inv[0:5]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size7 mux_bottom_track_1 (
		.in({chanx_right_in[33], chanx_right_in[69], chanx_right_in[103], chanx_left_in[1], chanx_left_in[7], chanx_left_in[37], chanx_left_in[73]}),
		.sram(mux_2level_tapbuf_size7_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_8_sram_inv[0:5]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size7 mux_bottom_track_9 (
		.in({chanx_right_in[32], chanx_right_in[68], chanx_right_in[99], chanx_left_in[2], chanx_left_in[11], chanx_left_in[38], chanx_left_in[74]}),
		.sram(mux_2level_tapbuf_size7_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_9_sram_inv[0:5]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size7 mux_bottom_track_185 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[38], chanx_right_in[74], chanx_left_in[32], chanx_left_in[68], chanx_left_in[99]}),
		.sram(mux_2level_tapbuf_size7_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_10_sram_inv[0:5]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size7 mux_bottom_track_193 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[37], chanx_right_in[73], chanx_left_in[33], chanx_left_in[69], chanx_left_in[103]}),
		.sram(mux_2level_tapbuf_size7_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_11_sram_inv[0:5]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size7 mux_bottom_track_201 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[36], chanx_right_in[72], chanx_left_in[34], chanx_left_in[70], chanx_left_in[104]}),
		.sram(mux_2level_tapbuf_size7_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_12_sram_inv[0:5]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size7 mux_bottom_track_209 (
		.in({chanx_right_in[34], chanx_right_in[70], chanx_right_in[104], chanx_left_in[0], chanx_left_in[3], chanx_left_in[36], chanx_left_in[72]}),
		.sram(mux_2level_tapbuf_size7_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_13_sram_inv[0:5]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size7 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[36], chany_top_in[72], chany_bottom_in[34], chany_bottom_in[70], chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size7_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_14_sram_inv[0:5]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size7 mux_left_track_9 (
		.in({chany_top_in[34], chany_top_in[70], chany_top_in[104], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[36], chany_bottom_in[72]}),
		.sram(mux_2level_tapbuf_size7_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_15_sram_inv[0:5]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size7 mux_left_track_17 (
		.in({chany_top_in[33], chany_top_in[69], chany_top_in[103], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size7_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_16_sram_inv[0:5]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size7 mux_left_track_25 (
		.in({chany_top_in[32], chany_top_in[68], chany_top_in[99], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[38], chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size7_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_17_sram_inv[0:5]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size7 mux_left_track_201 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[38], chany_top_in[74], chany_bottom_in[32], chany_bottom_in[68], chany_bottom_in[99]}),
		.sram(mux_2level_tapbuf_size7_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_18_sram_inv[0:5]),
		.out(chanx_left_out[100]));

	mux_2level_tapbuf_size7 mux_left_track_209 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[37], chany_top_in[73], chany_bottom_in[33], chany_bottom_in[69], chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size7_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_19_sram_inv[0:5]),
		.out(chanx_left_out[104]));

	mux_2level_tapbuf_size7_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_4_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_5_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_6_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_7_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_8_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_9_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_10_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_11_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_12_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_13_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_14_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_15_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_16_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_17_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_18_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_left_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_18_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_19_sram_inv[0:5]));

	mux_2level_tapbuf_size6 mux_right_track_0 (
		.in({chany_top_in[34], chany_top_in[70], chany_top_in[104], chany_bottom_in[33], chany_bottom_in[69], chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size6_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_0_sram_inv[0:5]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size6 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[69], chany_top_in[103], chany_bottom_in[34], chany_bottom_in[70], chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size6_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_1_sram_inv[0:5]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size6_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_0_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_1_sram_inv[0:5]));

endmodule
// ----- END Verilog module for sb_1__5_ -----

//----- Default net type -----
`default_nettype wire



