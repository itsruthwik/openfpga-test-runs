//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Sep 25 16:03:58 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__0_ -----
module sb_0__0_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:228] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:228] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:228] chany_top_out;
//----- OUTPUT PORTS -----
output [0:228] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_100_sram;
wire [0:1] mux_2level_tapbuf_size2_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_101_sram;
wire [0:1] mux_2level_tapbuf_size2_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_102_sram;
wire [0:1] mux_2level_tapbuf_size2_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_103_sram;
wire [0:1] mux_2level_tapbuf_size2_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_104_sram;
wire [0:1] mux_2level_tapbuf_size2_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_105_sram;
wire [0:1] mux_2level_tapbuf_size2_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_106_sram;
wire [0:1] mux_2level_tapbuf_size2_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_107_sram;
wire [0:1] mux_2level_tapbuf_size2_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_108_sram;
wire [0:1] mux_2level_tapbuf_size2_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_109_sram;
wire [0:1] mux_2level_tapbuf_size2_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_110_sram;
wire [0:1] mux_2level_tapbuf_size2_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_111_sram;
wire [0:1] mux_2level_tapbuf_size2_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_112_sram;
wire [0:1] mux_2level_tapbuf_size2_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_113_sram;
wire [0:1] mux_2level_tapbuf_size2_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_114_sram;
wire [0:1] mux_2level_tapbuf_size2_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_115_sram;
wire [0:1] mux_2level_tapbuf_size2_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_116_sram;
wire [0:1] mux_2level_tapbuf_size2_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_117_sram;
wire [0:1] mux_2level_tapbuf_size2_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_118_sram;
wire [0:1] mux_2level_tapbuf_size2_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_119_sram;
wire [0:1] mux_2level_tapbuf_size2_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_120_sram;
wire [0:1] mux_2level_tapbuf_size2_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_121_sram;
wire [0:1] mux_2level_tapbuf_size2_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_122_sram;
wire [0:1] mux_2level_tapbuf_size2_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_123_sram;
wire [0:1] mux_2level_tapbuf_size2_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_124_sram;
wire [0:1] mux_2level_tapbuf_size2_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_125_sram;
wire [0:1] mux_2level_tapbuf_size2_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_126_sram;
wire [0:1] mux_2level_tapbuf_size2_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_127_sram;
wire [0:1] mux_2level_tapbuf_size2_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_128_sram;
wire [0:1] mux_2level_tapbuf_size2_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_129_sram;
wire [0:1] mux_2level_tapbuf_size2_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_130_sram;
wire [0:1] mux_2level_tapbuf_size2_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_131_sram;
wire [0:1] mux_2level_tapbuf_size2_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_132_sram;
wire [0:1] mux_2level_tapbuf_size2_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_133_sram;
wire [0:1] mux_2level_tapbuf_size2_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_134_sram;
wire [0:1] mux_2level_tapbuf_size2_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_135_sram;
wire [0:1] mux_2level_tapbuf_size2_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_136_sram;
wire [0:1] mux_2level_tapbuf_size2_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_137_sram;
wire [0:1] mux_2level_tapbuf_size2_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_138_sram;
wire [0:1] mux_2level_tapbuf_size2_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_139_sram;
wire [0:1] mux_2level_tapbuf_size2_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_140_sram;
wire [0:1] mux_2level_tapbuf_size2_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_141_sram;
wire [0:1] mux_2level_tapbuf_size2_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_142_sram;
wire [0:1] mux_2level_tapbuf_size2_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_143_sram;
wire [0:1] mux_2level_tapbuf_size2_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_144_sram;
wire [0:1] mux_2level_tapbuf_size2_144_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_145_sram;
wire [0:1] mux_2level_tapbuf_size2_145_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_146_sram;
wire [0:1] mux_2level_tapbuf_size2_146_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_147_sram;
wire [0:1] mux_2level_tapbuf_size2_147_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_148_sram;
wire [0:1] mux_2level_tapbuf_size2_148_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_149_sram;
wire [0:1] mux_2level_tapbuf_size2_149_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_150_sram;
wire [0:1] mux_2level_tapbuf_size2_150_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_151_sram;
wire [0:1] mux_2level_tapbuf_size2_151_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_152_sram;
wire [0:1] mux_2level_tapbuf_size2_152_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_153_sram;
wire [0:1] mux_2level_tapbuf_size2_153_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_154_sram;
wire [0:1] mux_2level_tapbuf_size2_154_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_155_sram;
wire [0:1] mux_2level_tapbuf_size2_155_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_156_sram;
wire [0:1] mux_2level_tapbuf_size2_156_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_157_sram;
wire [0:1] mux_2level_tapbuf_size2_157_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_158_sram;
wire [0:1] mux_2level_tapbuf_size2_158_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_159_sram;
wire [0:1] mux_2level_tapbuf_size2_159_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_160_sram;
wire [0:1] mux_2level_tapbuf_size2_160_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_161_sram;
wire [0:1] mux_2level_tapbuf_size2_161_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_162_sram;
wire [0:1] mux_2level_tapbuf_size2_162_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_163_sram;
wire [0:1] mux_2level_tapbuf_size2_163_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_164_sram;
wire [0:1] mux_2level_tapbuf_size2_164_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_165_sram;
wire [0:1] mux_2level_tapbuf_size2_165_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_166_sram;
wire [0:1] mux_2level_tapbuf_size2_166_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_167_sram;
wire [0:1] mux_2level_tapbuf_size2_167_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_168_sram;
wire [0:1] mux_2level_tapbuf_size2_168_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_169_sram;
wire [0:1] mux_2level_tapbuf_size2_169_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_170_sram;
wire [0:1] mux_2level_tapbuf_size2_170_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_171_sram;
wire [0:1] mux_2level_tapbuf_size2_171_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_172_sram;
wire [0:1] mux_2level_tapbuf_size2_172_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_173_sram;
wire [0:1] mux_2level_tapbuf_size2_173_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_174_sram;
wire [0:1] mux_2level_tapbuf_size2_174_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_175_sram;
wire [0:1] mux_2level_tapbuf_size2_175_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_176_sram;
wire [0:1] mux_2level_tapbuf_size2_176_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_177_sram;
wire [0:1] mux_2level_tapbuf_size2_177_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_178_sram;
wire [0:1] mux_2level_tapbuf_size2_178_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_179_sram;
wire [0:1] mux_2level_tapbuf_size2_179_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_180_sram;
wire [0:1] mux_2level_tapbuf_size2_180_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_181_sram;
wire [0:1] mux_2level_tapbuf_size2_181_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_182_sram;
wire [0:1] mux_2level_tapbuf_size2_182_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_183_sram;
wire [0:1] mux_2level_tapbuf_size2_183_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_184_sram;
wire [0:1] mux_2level_tapbuf_size2_184_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_185_sram;
wire [0:1] mux_2level_tapbuf_size2_185_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_186_sram;
wire [0:1] mux_2level_tapbuf_size2_186_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_187_sram;
wire [0:1] mux_2level_tapbuf_size2_187_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_188_sram;
wire [0:1] mux_2level_tapbuf_size2_188_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_189_sram;
wire [0:1] mux_2level_tapbuf_size2_189_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_190_sram;
wire [0:1] mux_2level_tapbuf_size2_190_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_191_sram;
wire [0:1] mux_2level_tapbuf_size2_191_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_192_sram;
wire [0:1] mux_2level_tapbuf_size2_192_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_193_sram;
wire [0:1] mux_2level_tapbuf_size2_193_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_194_sram;
wire [0:1] mux_2level_tapbuf_size2_194_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_195_sram;
wire [0:1] mux_2level_tapbuf_size2_195_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_196_sram;
wire [0:1] mux_2level_tapbuf_size2_196_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_197_sram;
wire [0:1] mux_2level_tapbuf_size2_197_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_198_sram;
wire [0:1] mux_2level_tapbuf_size2_198_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_199_sram;
wire [0:1] mux_2level_tapbuf_size2_199_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_200_sram;
wire [0:1] mux_2level_tapbuf_size2_200_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_201_sram;
wire [0:1] mux_2level_tapbuf_size2_201_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_202_sram;
wire [0:1] mux_2level_tapbuf_size2_202_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_203_sram;
wire [0:1] mux_2level_tapbuf_size2_203_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_204_sram;
wire [0:1] mux_2level_tapbuf_size2_204_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_205_sram;
wire [0:1] mux_2level_tapbuf_size2_205_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_206_sram;
wire [0:1] mux_2level_tapbuf_size2_206_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_207_sram;
wire [0:1] mux_2level_tapbuf_size2_207_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_208_sram;
wire [0:1] mux_2level_tapbuf_size2_208_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_209_sram;
wire [0:1] mux_2level_tapbuf_size2_209_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_210_sram;
wire [0:1] mux_2level_tapbuf_size2_210_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_211_sram;
wire [0:1] mux_2level_tapbuf_size2_211_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_212_sram;
wire [0:1] mux_2level_tapbuf_size2_212_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_213_sram;
wire [0:1] mux_2level_tapbuf_size2_213_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_214_sram;
wire [0:1] mux_2level_tapbuf_size2_214_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_215_sram;
wire [0:1] mux_2level_tapbuf_size2_215_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_216_sram;
wire [0:1] mux_2level_tapbuf_size2_216_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_217_sram;
wire [0:1] mux_2level_tapbuf_size2_217_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_218_sram;
wire [0:1] mux_2level_tapbuf_size2_218_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_219_sram;
wire [0:1] mux_2level_tapbuf_size2_219_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_220_sram;
wire [0:1] mux_2level_tapbuf_size2_220_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_221_sram;
wire [0:1] mux_2level_tapbuf_size2_221_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_222_sram;
wire [0:1] mux_2level_tapbuf_size2_222_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_223_sram;
wire [0:1] mux_2level_tapbuf_size2_223_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_224_sram;
wire [0:1] mux_2level_tapbuf_size2_224_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_225_sram;
wire [0:1] mux_2level_tapbuf_size2_225_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_226_sram;
wire [0:1] mux_2level_tapbuf_size2_226_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_227_sram;
wire [0:1] mux_2level_tapbuf_size2_227_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_228_sram;
wire [0:1] mux_2level_tapbuf_size2_228_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_229_sram;
wire [0:1] mux_2level_tapbuf_size2_229_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_230_sram;
wire [0:1] mux_2level_tapbuf_size2_230_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_231_sram;
wire [0:1] mux_2level_tapbuf_size2_231_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_232_sram;
wire [0:1] mux_2level_tapbuf_size2_232_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_233_sram;
wire [0:1] mux_2level_tapbuf_size2_233_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_234_sram;
wire [0:1] mux_2level_tapbuf_size2_234_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_235_sram;
wire [0:1] mux_2level_tapbuf_size2_235_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_236_sram;
wire [0:1] mux_2level_tapbuf_size2_236_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_237_sram;
wire [0:1] mux_2level_tapbuf_size2_237_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_238_sram;
wire [0:1] mux_2level_tapbuf_size2_238_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_239_sram;
wire [0:1] mux_2level_tapbuf_size2_239_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_240_sram;
wire [0:1] mux_2level_tapbuf_size2_240_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_241_sram;
wire [0:1] mux_2level_tapbuf_size2_241_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_242_sram;
wire [0:1] mux_2level_tapbuf_size2_242_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_243_sram;
wire [0:1] mux_2level_tapbuf_size2_243_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_244_sram;
wire [0:1] mux_2level_tapbuf_size2_244_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_245_sram;
wire [0:1] mux_2level_tapbuf_size2_245_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_246_sram;
wire [0:1] mux_2level_tapbuf_size2_246_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_247_sram;
wire [0:1] mux_2level_tapbuf_size2_247_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_248_sram;
wire [0:1] mux_2level_tapbuf_size2_248_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_249_sram;
wire [0:1] mux_2level_tapbuf_size2_249_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_250_sram;
wire [0:1] mux_2level_tapbuf_size2_250_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_251_sram;
wire [0:1] mux_2level_tapbuf_size2_251_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_252_sram;
wire [0:1] mux_2level_tapbuf_size2_252_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_253_sram;
wire [0:1] mux_2level_tapbuf_size2_253_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_254_sram;
wire [0:1] mux_2level_tapbuf_size2_254_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_255_sram;
wire [0:1] mux_2level_tapbuf_size2_255_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_256_sram;
wire [0:1] mux_2level_tapbuf_size2_256_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_257_sram;
wire [0:1] mux_2level_tapbuf_size2_257_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_258_sram;
wire [0:1] mux_2level_tapbuf_size2_258_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_259_sram;
wire [0:1] mux_2level_tapbuf_size2_259_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_260_sram;
wire [0:1] mux_2level_tapbuf_size2_260_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_261_sram;
wire [0:1] mux_2level_tapbuf_size2_261_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_262_sram;
wire [0:1] mux_2level_tapbuf_size2_262_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_263_sram;
wire [0:1] mux_2level_tapbuf_size2_263_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_264_sram;
wire [0:1] mux_2level_tapbuf_size2_264_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_265_sram;
wire [0:1] mux_2level_tapbuf_size2_265_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_266_sram;
wire [0:1] mux_2level_tapbuf_size2_266_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_267_sram;
wire [0:1] mux_2level_tapbuf_size2_267_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_268_sram;
wire [0:1] mux_2level_tapbuf_size2_268_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_269_sram;
wire [0:1] mux_2level_tapbuf_size2_269_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_270_sram;
wire [0:1] mux_2level_tapbuf_size2_270_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_271_sram;
wire [0:1] mux_2level_tapbuf_size2_271_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_272_sram;
wire [0:1] mux_2level_tapbuf_size2_272_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_273_sram;
wire [0:1] mux_2level_tapbuf_size2_273_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_274_sram;
wire [0:1] mux_2level_tapbuf_size2_274_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_275_sram;
wire [0:1] mux_2level_tapbuf_size2_275_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_276_sram;
wire [0:1] mux_2level_tapbuf_size2_276_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_277_sram;
wire [0:1] mux_2level_tapbuf_size2_277_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_278_sram;
wire [0:1] mux_2level_tapbuf_size2_278_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_279_sram;
wire [0:1] mux_2level_tapbuf_size2_279_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_280_sram;
wire [0:1] mux_2level_tapbuf_size2_280_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_281_sram;
wire [0:1] mux_2level_tapbuf_size2_281_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_282_sram;
wire [0:1] mux_2level_tapbuf_size2_282_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_283_sram;
wire [0:1] mux_2level_tapbuf_size2_283_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_284_sram;
wire [0:1] mux_2level_tapbuf_size2_284_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_285_sram;
wire [0:1] mux_2level_tapbuf_size2_285_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_286_sram;
wire [0:1] mux_2level_tapbuf_size2_286_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_287_sram;
wire [0:1] mux_2level_tapbuf_size2_287_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_288_sram;
wire [0:1] mux_2level_tapbuf_size2_288_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_289_sram;
wire [0:1] mux_2level_tapbuf_size2_289_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_290_sram;
wire [0:1] mux_2level_tapbuf_size2_290_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_291_sram;
wire [0:1] mux_2level_tapbuf_size2_291_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_292_sram;
wire [0:1] mux_2level_tapbuf_size2_292_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_293_sram;
wire [0:1] mux_2level_tapbuf_size2_293_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_294_sram;
wire [0:1] mux_2level_tapbuf_size2_294_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_295_sram;
wire [0:1] mux_2level_tapbuf_size2_295_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_296_sram;
wire [0:1] mux_2level_tapbuf_size2_296_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_297_sram;
wire [0:1] mux_2level_tapbuf_size2_297_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_298_sram;
wire [0:1] mux_2level_tapbuf_size2_298_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_299_sram;
wire [0:1] mux_2level_tapbuf_size2_299_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_300_sram;
wire [0:1] mux_2level_tapbuf_size2_300_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_301_sram;
wire [0:1] mux_2level_tapbuf_size2_301_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_302_sram;
wire [0:1] mux_2level_tapbuf_size2_302_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_303_sram;
wire [0:1] mux_2level_tapbuf_size2_303_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_304_sram;
wire [0:1] mux_2level_tapbuf_size2_304_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_305_sram;
wire [0:1] mux_2level_tapbuf_size2_305_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_306_sram;
wire [0:1] mux_2level_tapbuf_size2_306_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_307_sram;
wire [0:1] mux_2level_tapbuf_size2_307_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_308_sram;
wire [0:1] mux_2level_tapbuf_size2_308_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_309_sram;
wire [0:1] mux_2level_tapbuf_size2_309_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_310_sram;
wire [0:1] mux_2level_tapbuf_size2_310_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_311_sram;
wire [0:1] mux_2level_tapbuf_size2_311_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_312_sram;
wire [0:1] mux_2level_tapbuf_size2_312_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_313_sram;
wire [0:1] mux_2level_tapbuf_size2_313_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_314_sram;
wire [0:1] mux_2level_tapbuf_size2_314_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_315_sram;
wire [0:1] mux_2level_tapbuf_size2_315_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_316_sram;
wire [0:1] mux_2level_tapbuf_size2_316_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_317_sram;
wire [0:1] mux_2level_tapbuf_size2_317_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_318_sram;
wire [0:1] mux_2level_tapbuf_size2_318_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_319_sram;
wire [0:1] mux_2level_tapbuf_size2_319_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_320_sram;
wire [0:1] mux_2level_tapbuf_size2_320_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_321_sram;
wire [0:1] mux_2level_tapbuf_size2_321_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_322_sram;
wire [0:1] mux_2level_tapbuf_size2_322_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_323_sram;
wire [0:1] mux_2level_tapbuf_size2_323_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_324_sram;
wire [0:1] mux_2level_tapbuf_size2_324_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_325_sram;
wire [0:1] mux_2level_tapbuf_size2_325_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_326_sram;
wire [0:1] mux_2level_tapbuf_size2_326_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_327_sram;
wire [0:1] mux_2level_tapbuf_size2_327_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_328_sram;
wire [0:1] mux_2level_tapbuf_size2_328_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_329_sram;
wire [0:1] mux_2level_tapbuf_size2_329_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_330_sram;
wire [0:1] mux_2level_tapbuf_size2_330_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_331_sram;
wire [0:1] mux_2level_tapbuf_size2_331_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_332_sram;
wire [0:1] mux_2level_tapbuf_size2_332_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_333_sram;
wire [0:1] mux_2level_tapbuf_size2_333_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_334_sram;
wire [0:1] mux_2level_tapbuf_size2_334_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_335_sram;
wire [0:1] mux_2level_tapbuf_size2_335_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_336_sram;
wire [0:1] mux_2level_tapbuf_size2_336_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_337_sram;
wire [0:1] mux_2level_tapbuf_size2_337_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_338_sram;
wire [0:1] mux_2level_tapbuf_size2_338_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_339_sram;
wire [0:1] mux_2level_tapbuf_size2_339_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_340_sram;
wire [0:1] mux_2level_tapbuf_size2_340_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_341_sram;
wire [0:1] mux_2level_tapbuf_size2_341_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_342_sram;
wire [0:1] mux_2level_tapbuf_size2_342_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_343_sram;
wire [0:1] mux_2level_tapbuf_size2_343_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_344_sram;
wire [0:1] mux_2level_tapbuf_size2_344_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_345_sram;
wire [0:1] mux_2level_tapbuf_size2_345_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_346_sram;
wire [0:1] mux_2level_tapbuf_size2_346_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_347_sram;
wire [0:1] mux_2level_tapbuf_size2_347_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_348_sram;
wire [0:1] mux_2level_tapbuf_size2_348_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_349_sram;
wire [0:1] mux_2level_tapbuf_size2_349_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_350_sram;
wire [0:1] mux_2level_tapbuf_size2_350_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_351_sram;
wire [0:1] mux_2level_tapbuf_size2_351_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_352_sram;
wire [0:1] mux_2level_tapbuf_size2_352_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_353_sram;
wire [0:1] mux_2level_tapbuf_size2_353_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_354_sram;
wire [0:1] mux_2level_tapbuf_size2_354_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_355_sram;
wire [0:1] mux_2level_tapbuf_size2_355_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_356_sram;
wire [0:1] mux_2level_tapbuf_size2_356_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_357_sram;
wire [0:1] mux_2level_tapbuf_size2_357_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_358_sram;
wire [0:1] mux_2level_tapbuf_size2_358_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_359_sram;
wire [0:1] mux_2level_tapbuf_size2_359_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_360_sram;
wire [0:1] mux_2level_tapbuf_size2_360_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_361_sram;
wire [0:1] mux_2level_tapbuf_size2_361_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_362_sram;
wire [0:1] mux_2level_tapbuf_size2_362_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_363_sram;
wire [0:1] mux_2level_tapbuf_size2_363_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_364_sram;
wire [0:1] mux_2level_tapbuf_size2_364_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_365_sram;
wire [0:1] mux_2level_tapbuf_size2_365_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_366_sram;
wire [0:1] mux_2level_tapbuf_size2_366_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_367_sram;
wire [0:1] mux_2level_tapbuf_size2_367_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_368_sram;
wire [0:1] mux_2level_tapbuf_size2_368_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_369_sram;
wire [0:1] mux_2level_tapbuf_size2_369_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_370_sram;
wire [0:1] mux_2level_tapbuf_size2_370_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_371_sram;
wire [0:1] mux_2level_tapbuf_size2_371_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_372_sram;
wire [0:1] mux_2level_tapbuf_size2_372_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_373_sram;
wire [0:1] mux_2level_tapbuf_size2_373_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_374_sram;
wire [0:1] mux_2level_tapbuf_size2_374_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_375_sram;
wire [0:1] mux_2level_tapbuf_size2_375_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_376_sram;
wire [0:1] mux_2level_tapbuf_size2_376_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_377_sram;
wire [0:1] mux_2level_tapbuf_size2_377_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_378_sram;
wire [0:1] mux_2level_tapbuf_size2_378_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_379_sram;
wire [0:1] mux_2level_tapbuf_size2_379_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_380_sram;
wire [0:1] mux_2level_tapbuf_size2_380_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_381_sram;
wire [0:1] mux_2level_tapbuf_size2_381_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_382_sram;
wire [0:1] mux_2level_tapbuf_size2_382_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_383_sram;
wire [0:1] mux_2level_tapbuf_size2_383_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_384_sram;
wire [0:1] mux_2level_tapbuf_size2_384_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_385_sram;
wire [0:1] mux_2level_tapbuf_size2_385_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_386_sram;
wire [0:1] mux_2level_tapbuf_size2_386_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_387_sram;
wire [0:1] mux_2level_tapbuf_size2_387_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_388_sram;
wire [0:1] mux_2level_tapbuf_size2_388_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_389_sram;
wire [0:1] mux_2level_tapbuf_size2_389_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_390_sram;
wire [0:1] mux_2level_tapbuf_size2_390_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_391_sram;
wire [0:1] mux_2level_tapbuf_size2_391_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_392_sram;
wire [0:1] mux_2level_tapbuf_size2_392_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_393_sram;
wire [0:1] mux_2level_tapbuf_size2_393_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_394_sram;
wire [0:1] mux_2level_tapbuf_size2_394_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_395_sram;
wire [0:1] mux_2level_tapbuf_size2_395_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_396_sram;
wire [0:1] mux_2level_tapbuf_size2_396_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_397_sram;
wire [0:1] mux_2level_tapbuf_size2_397_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_398_sram;
wire [0:1] mux_2level_tapbuf_size2_398_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_399_sram;
wire [0:1] mux_2level_tapbuf_size2_399_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_60_sram;
wire [0:1] mux_2level_tapbuf_size2_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_61_sram;
wire [0:1] mux_2level_tapbuf_size2_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_62_sram;
wire [0:1] mux_2level_tapbuf_size2_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_63_sram;
wire [0:1] mux_2level_tapbuf_size2_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_64_sram;
wire [0:1] mux_2level_tapbuf_size2_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_65_sram;
wire [0:1] mux_2level_tapbuf_size2_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_66_sram;
wire [0:1] mux_2level_tapbuf_size2_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_67_sram;
wire [0:1] mux_2level_tapbuf_size2_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_68_sram;
wire [0:1] mux_2level_tapbuf_size2_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_69_sram;
wire [0:1] mux_2level_tapbuf_size2_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_70_sram;
wire [0:1] mux_2level_tapbuf_size2_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_71_sram;
wire [0:1] mux_2level_tapbuf_size2_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_72_sram;
wire [0:1] mux_2level_tapbuf_size2_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_73_sram;
wire [0:1] mux_2level_tapbuf_size2_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_74_sram;
wire [0:1] mux_2level_tapbuf_size2_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_75_sram;
wire [0:1] mux_2level_tapbuf_size2_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_76_sram;
wire [0:1] mux_2level_tapbuf_size2_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_77_sram;
wire [0:1] mux_2level_tapbuf_size2_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_78_sram;
wire [0:1] mux_2level_tapbuf_size2_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_79_sram;
wire [0:1] mux_2level_tapbuf_size2_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_80_sram;
wire [0:1] mux_2level_tapbuf_size2_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_81_sram;
wire [0:1] mux_2level_tapbuf_size2_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_82_sram;
wire [0:1] mux_2level_tapbuf_size2_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_83_sram;
wire [0:1] mux_2level_tapbuf_size2_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_84_sram;
wire [0:1] mux_2level_tapbuf_size2_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_85_sram;
wire [0:1] mux_2level_tapbuf_size2_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_86_sram;
wire [0:1] mux_2level_tapbuf_size2_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_87_sram;
wire [0:1] mux_2level_tapbuf_size2_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_88_sram;
wire [0:1] mux_2level_tapbuf_size2_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_89_sram;
wire [0:1] mux_2level_tapbuf_size2_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_90_sram;
wire [0:1] mux_2level_tapbuf_size2_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_91_sram;
wire [0:1] mux_2level_tapbuf_size2_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_92_sram;
wire [0:1] mux_2level_tapbuf_size2_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_93_sram;
wire [0:1] mux_2level_tapbuf_size2_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_94_sram;
wire [0:1] mux_2level_tapbuf_size2_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_95_sram;
wire [0:1] mux_2level_tapbuf_size2_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_96_sram;
wire [0:1] mux_2level_tapbuf_size2_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_97_sram;
wire [0:1] mux_2level_tapbuf_size2_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_98_sram;
wire [0:1] mux_2level_tapbuf_size2_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_99_sram;
wire [0:1] mux_2level_tapbuf_size2_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_144_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_145_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_146_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_147_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_148_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_149_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_150_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_151_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_152_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_153_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_154_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_155_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_156_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_157_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_158_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_159_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_160_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_161_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_162_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_163_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_164_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_165_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_166_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_167_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_168_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_169_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_170_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_171_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_172_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_173_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_174_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_175_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_176_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_177_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_178_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_179_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_180_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_181_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_182_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_183_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_184_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_185_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_186_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_187_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_188_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_189_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_190_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_191_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_192_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_193_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_194_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_195_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_196_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_197_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_198_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_199_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_200_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_201_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_202_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_203_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_204_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_205_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_206_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_207_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_208_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_209_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_210_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_211_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_212_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_213_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_214_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_215_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_216_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_217_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_218_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_219_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_220_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_221_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_222_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_223_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_224_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_225_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_226_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_227_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_228_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_229_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_230_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_231_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_232_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_233_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_234_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_235_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_236_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_237_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_238_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_239_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_240_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_241_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_242_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_243_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_244_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_245_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_246_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_247_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_248_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_249_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_250_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_251_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_252_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_253_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_254_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_255_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_256_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_257_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_258_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_259_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_260_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_261_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_262_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_263_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_264_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_265_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_266_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_267_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_268_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_269_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_270_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_271_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_272_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_273_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_274_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_275_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_276_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_277_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_278_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_279_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_280_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_281_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_282_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_283_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_284_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_285_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_286_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_287_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_288_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_289_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_290_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_291_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_292_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_293_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_294_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_295_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_296_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_297_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_298_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_299_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_300_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_301_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_302_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_303_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_304_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_305_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_306_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_307_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_308_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_309_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_310_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_311_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_312_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_313_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_314_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_315_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_316_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_317_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_318_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_319_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_320_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_321_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_322_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_323_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_324_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_325_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_326_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_327_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_328_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_329_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_330_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_331_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_332_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_333_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_334_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_335_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_336_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_337_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_338_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_339_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_340_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_341_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_342_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_343_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_344_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_345_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_346_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_347_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_348_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_349_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_350_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_351_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_352_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_353_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_354_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_355_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_356_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_357_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_358_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_359_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_360_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_361_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_362_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_363_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_364_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_365_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_366_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_367_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_368_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_369_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_370_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_371_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_372_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_373_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_374_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_375_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_376_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_377_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_378_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_379_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_380_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_381_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_382_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_383_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_384_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_385_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_386_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_387_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_388_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_389_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_390_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_391_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_392_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_393_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_394_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_395_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_396_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_397_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_398_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chany_top_in[7];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chany_top_in[43];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[80] = chany_top_in[79];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[116] = chany_top_in[115];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[152] = chany_top_in[151];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[188] = chany_top_in[187];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[197] = chany_top_in[196];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[206] = chany_top_in[205];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[215] = chany_top_in[214];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[224] = chany_top_in[223];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chanx_right_in[9];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chanx_right_in[18];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chanx_right_in[27];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chanx_right_in[36];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chanx_right_in[45];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chanx_right_in[54];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chanx_right_in[63];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chanx_right_in[72];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chanx_right_in[81];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chanx_right_in[90];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chanx_right_in[99];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chanx_right_in[108];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chanx_right_in[117];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chanx_right_in[126];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chanx_right_in[135];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chanx_right_in[144];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chanx_right_in[153];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chanx_right_in[162];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chanx_right_in[171];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chanx_right_in[180];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[188] = chanx_right_in[189];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chanx_right_in[198];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chanx_right_in[207];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chanx_right_in[216];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[224] = chanx_right_in[225];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size3 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[1]}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size3 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[2]}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_2level_tapbuf_size3 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[3]}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size3 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[4]}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_2level_tapbuf_size3 mux_right_track_0 (
		.in({chany_top_in[228], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[0], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size3_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_199_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[5]}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size2 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[6]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_2level_tapbuf_size2 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[7]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size2 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[8]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_2level_tapbuf_size2 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[10]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_2level_tapbuf_size2 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[11]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size2 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[12]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_2level_tapbuf_size2 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[13]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size2 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[14]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_2level_tapbuf_size2 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[15]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size2 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[16]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_2level_tapbuf_size2 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[17]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size2 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[19]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size2 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[20]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_2level_tapbuf_size2 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[21]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size2 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[22]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_2level_tapbuf_size2 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[23]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size2 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[24]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_2level_tapbuf_size2 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[25]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size2 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[26]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_2level_tapbuf_size2 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[28]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_2level_tapbuf_size2 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[29]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size2 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[30]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_2level_tapbuf_size2 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[31]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size2 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[32]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_2level_tapbuf_size2 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[33]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size2 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[34]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_2level_tapbuf_size2 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[35]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size2 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[37]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size2 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[38]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_2level_tapbuf_size2 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[39]}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size2 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[40]}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_2level_tapbuf_size2 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[41]}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size2 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[42]}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_2level_tapbuf_size2 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[43]}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size2 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[44]}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_2level_tapbuf_size2 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[46]}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_2level_tapbuf_size2 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[47]}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size2 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[48]}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_2level_tapbuf_size2 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[49]}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size2 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[50]}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_2level_tapbuf_size2 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[51]}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size2 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[52]}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_2level_tapbuf_size2 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[53]}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size2 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[55]}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size2 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[56]}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_2level_tapbuf_size2 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[57]}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size2 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[58]}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_2level_tapbuf_size2 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[59]}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size2 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[60]}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_2level_tapbuf_size2 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[61]}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size2 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[62]}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_2level_tapbuf_size2 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[64]}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_2level_tapbuf_size2 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[65]}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size2 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[66]}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_2level_tapbuf_size2 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[67]}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size2 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[68]}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_2level_tapbuf_size2 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[69]}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size2 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[70]}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_2level_tapbuf_size2 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[71]}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size2 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[73]}),
		.sram(mux_2level_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_60_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size2 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[74]}),
		.sram(mux_2level_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_61_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_2level_tapbuf_size2 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[75]}),
		.sram(mux_2level_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_62_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size2 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[76]}),
		.sram(mux_2level_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_63_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_2level_tapbuf_size2 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[77]}),
		.sram(mux_2level_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_64_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size2 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[78]}),
		.sram(mux_2level_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_65_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_2level_tapbuf_size2 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[79]}),
		.sram(mux_2level_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_66_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size2 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[80]}),
		.sram(mux_2level_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_67_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_2level_tapbuf_size2 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[82]}),
		.sram(mux_2level_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_68_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_2level_tapbuf_size2 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[83]}),
		.sram(mux_2level_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_69_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size2 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[84]}),
		.sram(mux_2level_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_70_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_2level_tapbuf_size2 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[85]}),
		.sram(mux_2level_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_71_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size2 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[86]}),
		.sram(mux_2level_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_72_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_2level_tapbuf_size2 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[87]}),
		.sram(mux_2level_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_73_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size2 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[88]}),
		.sram(mux_2level_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_74_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_2level_tapbuf_size2 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[89]}),
		.sram(mux_2level_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_75_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size2 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[91]}),
		.sram(mux_2level_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_76_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size2 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[92]}),
		.sram(mux_2level_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_77_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_2level_tapbuf_size2 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[93]}),
		.sram(mux_2level_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_78_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size2 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[94]}),
		.sram(mux_2level_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_79_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_2level_tapbuf_size2 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[95]}),
		.sram(mux_2level_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_80_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size2 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[96]}),
		.sram(mux_2level_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_81_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_2level_tapbuf_size2 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[97]}),
		.sram(mux_2level_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_82_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size2 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[98]}),
		.sram(mux_2level_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_83_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_2level_tapbuf_size2 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[100]}),
		.sram(mux_2level_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_84_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_2level_tapbuf_size2 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[101]}),
		.sram(mux_2level_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_85_sram_inv[0:1]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size2 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[102]}),
		.sram(mux_2level_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_86_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_2level_tapbuf_size2 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[103]}),
		.sram(mux_2level_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_87_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size2 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[104]}),
		.sram(mux_2level_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_88_sram_inv[0:1]),
		.out(chany_top_out[103]));

	mux_2level_tapbuf_size2 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[105]}),
		.sram(mux_2level_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_89_sram_inv[0:1]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size2 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[106]}),
		.sram(mux_2level_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_90_sram_inv[0:1]),
		.out(chany_top_out[105]));

	mux_2level_tapbuf_size2 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[107]}),
		.sram(mux_2level_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_91_sram_inv[0:1]),
		.out(chany_top_out[106]));

	mux_2level_tapbuf_size2 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[109]}),
		.sram(mux_2level_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_92_sram_inv[0:1]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size2 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[110]}),
		.sram(mux_2level_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_93_sram_inv[0:1]),
		.out(chany_top_out[109]));

	mux_2level_tapbuf_size2 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[111]}),
		.sram(mux_2level_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_94_sram_inv[0:1]),
		.out(chany_top_out[110]));

	mux_2level_tapbuf_size2 mux_top_track_222 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[112]}),
		.sram(mux_2level_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_95_sram_inv[0:1]),
		.out(chany_top_out[111]));

	mux_2level_tapbuf_size2 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[113]}),
		.sram(mux_2level_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_96_sram_inv[0:1]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size2 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[114]}),
		.sram(mux_2level_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_97_sram_inv[0:1]),
		.out(chany_top_out[113]));

	mux_2level_tapbuf_size2 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[115]}),
		.sram(mux_2level_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_98_sram_inv[0:1]),
		.out(chany_top_out[114]));

	mux_2level_tapbuf_size2 mux_top_track_230 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[116]}),
		.sram(mux_2level_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_99_sram_inv[0:1]),
		.out(chany_top_out[115]));

	mux_2level_tapbuf_size2 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[118]}),
		.sram(mux_2level_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_100_sram_inv[0:1]),
		.out(chany_top_out[117]));

	mux_2level_tapbuf_size2 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[119]}),
		.sram(mux_2level_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_101_sram_inv[0:1]),
		.out(chany_top_out[118]));

	mux_2level_tapbuf_size2 mux_top_track_238 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[120]}),
		.sram(mux_2level_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_102_sram_inv[0:1]),
		.out(chany_top_out[119]));

	mux_2level_tapbuf_size2 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[121]}),
		.sram(mux_2level_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_103_sram_inv[0:1]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size2 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[122]}),
		.sram(mux_2level_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_104_sram_inv[0:1]),
		.out(chany_top_out[121]));

	mux_2level_tapbuf_size2 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[123]}),
		.sram(mux_2level_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_105_sram_inv[0:1]),
		.out(chany_top_out[122]));

	mux_2level_tapbuf_size2 mux_top_track_246 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[124]}),
		.sram(mux_2level_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_106_sram_inv[0:1]),
		.out(chany_top_out[123]));

	mux_2level_tapbuf_size2 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[125]}),
		.sram(mux_2level_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_107_sram_inv[0:1]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size2 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[127]}),
		.sram(mux_2level_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_108_sram_inv[0:1]),
		.out(chany_top_out[126]));

	mux_2level_tapbuf_size2 mux_top_track_254 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[128]}),
		.sram(mux_2level_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_109_sram_inv[0:1]),
		.out(chany_top_out[127]));

	mux_2level_tapbuf_size2 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[129]}),
		.sram(mux_2level_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_110_sram_inv[0:1]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size2 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[130]}),
		.sram(mux_2level_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_111_sram_inv[0:1]),
		.out(chany_top_out[129]));

	mux_2level_tapbuf_size2 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[131]}),
		.sram(mux_2level_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_112_sram_inv[0:1]),
		.out(chany_top_out[130]));

	mux_2level_tapbuf_size2 mux_top_track_262 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[132]}),
		.sram(mux_2level_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_113_sram_inv[0:1]),
		.out(chany_top_out[131]));

	mux_2level_tapbuf_size2 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[133]}),
		.sram(mux_2level_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_114_sram_inv[0:1]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size2 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[134]}),
		.sram(mux_2level_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_115_sram_inv[0:1]),
		.out(chany_top_out[133]));

	mux_2level_tapbuf_size2 mux_top_track_270 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[136]}),
		.sram(mux_2level_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_116_sram_inv[0:1]),
		.out(chany_top_out[135]));

	mux_2level_tapbuf_size2 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[137]}),
		.sram(mux_2level_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_117_sram_inv[0:1]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size2 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[138]}),
		.sram(mux_2level_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_118_sram_inv[0:1]),
		.out(chany_top_out[137]));

	mux_2level_tapbuf_size2 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[139]}),
		.sram(mux_2level_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_119_sram_inv[0:1]),
		.out(chany_top_out[138]));

	mux_2level_tapbuf_size2 mux_top_track_278 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[140]}),
		.sram(mux_2level_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_120_sram_inv[0:1]),
		.out(chany_top_out[139]));

	mux_2level_tapbuf_size2 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[141]}),
		.sram(mux_2level_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_121_sram_inv[0:1]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size2 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[142]}),
		.sram(mux_2level_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_122_sram_inv[0:1]),
		.out(chany_top_out[141]));

	mux_2level_tapbuf_size2 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[143]}),
		.sram(mux_2level_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_123_sram_inv[0:1]),
		.out(chany_top_out[142]));

	mux_2level_tapbuf_size2 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[145]}),
		.sram(mux_2level_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_124_sram_inv[0:1]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size2 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[146]}),
		.sram(mux_2level_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_125_sram_inv[0:1]),
		.out(chany_top_out[145]));

	mux_2level_tapbuf_size2 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[147]}),
		.sram(mux_2level_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_126_sram_inv[0:1]),
		.out(chany_top_out[146]));

	mux_2level_tapbuf_size2 mux_top_track_294 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[148]}),
		.sram(mux_2level_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_127_sram_inv[0:1]),
		.out(chany_top_out[147]));

	mux_2level_tapbuf_size2 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[149]}),
		.sram(mux_2level_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_128_sram_inv[0:1]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size2 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[150]}),
		.sram(mux_2level_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_129_sram_inv[0:1]),
		.out(chany_top_out[149]));

	mux_2level_tapbuf_size2 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[151]}),
		.sram(mux_2level_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_130_sram_inv[0:1]),
		.out(chany_top_out[150]));

	mux_2level_tapbuf_size2 mux_top_track_302 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[152]}),
		.sram(mux_2level_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_131_sram_inv[0:1]),
		.out(chany_top_out[151]));

	mux_2level_tapbuf_size2 mux_top_track_306 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[154]}),
		.sram(mux_2level_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_132_sram_inv[0:1]),
		.out(chany_top_out[153]));

	mux_2level_tapbuf_size2 mux_top_track_308 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[155]}),
		.sram(mux_2level_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_133_sram_inv[0:1]),
		.out(chany_top_out[154]));

	mux_2level_tapbuf_size2 mux_top_track_310 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[156]}),
		.sram(mux_2level_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_134_sram_inv[0:1]),
		.out(chany_top_out[155]));

	mux_2level_tapbuf_size2 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[157]}),
		.sram(mux_2level_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_135_sram_inv[0:1]),
		.out(chany_top_out[156]));

	mux_2level_tapbuf_size2 mux_top_track_314 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[158]}),
		.sram(mux_2level_tapbuf_size2_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_136_sram_inv[0:1]),
		.out(chany_top_out[157]));

	mux_2level_tapbuf_size2 mux_top_track_316 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[159]}),
		.sram(mux_2level_tapbuf_size2_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_137_sram_inv[0:1]),
		.out(chany_top_out[158]));

	mux_2level_tapbuf_size2 mux_top_track_318 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[160]}),
		.sram(mux_2level_tapbuf_size2_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_138_sram_inv[0:1]),
		.out(chany_top_out[159]));

	mux_2level_tapbuf_size2 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[161]}),
		.sram(mux_2level_tapbuf_size2_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_139_sram_inv[0:1]),
		.out(chany_top_out[160]));

	mux_2level_tapbuf_size2 mux_top_track_324 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[163]}),
		.sram(mux_2level_tapbuf_size2_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_140_sram_inv[0:1]),
		.out(chany_top_out[162]));

	mux_2level_tapbuf_size2 mux_top_track_326 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[164]}),
		.sram(mux_2level_tapbuf_size2_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_141_sram_inv[0:1]),
		.out(chany_top_out[163]));

	mux_2level_tapbuf_size2 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[165]}),
		.sram(mux_2level_tapbuf_size2_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_142_sram_inv[0:1]),
		.out(chany_top_out[164]));

	mux_2level_tapbuf_size2 mux_top_track_330 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[166]}),
		.sram(mux_2level_tapbuf_size2_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_143_sram_inv[0:1]),
		.out(chany_top_out[165]));

	mux_2level_tapbuf_size2 mux_top_track_332 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[167]}),
		.sram(mux_2level_tapbuf_size2_144_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_144_sram_inv[0:1]),
		.out(chany_top_out[166]));

	mux_2level_tapbuf_size2 mux_top_track_334 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[168]}),
		.sram(mux_2level_tapbuf_size2_145_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_145_sram_inv[0:1]),
		.out(chany_top_out[167]));

	mux_2level_tapbuf_size2 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[169]}),
		.sram(mux_2level_tapbuf_size2_146_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_146_sram_inv[0:1]),
		.out(chany_top_out[168]));

	mux_2level_tapbuf_size2 mux_top_track_338 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[170]}),
		.sram(mux_2level_tapbuf_size2_147_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_147_sram_inv[0:1]),
		.out(chany_top_out[169]));

	mux_2level_tapbuf_size2 mux_top_track_342 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[172]}),
		.sram(mux_2level_tapbuf_size2_148_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_148_sram_inv[0:1]),
		.out(chany_top_out[171]));

	mux_2level_tapbuf_size2 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[173]}),
		.sram(mux_2level_tapbuf_size2_149_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_149_sram_inv[0:1]),
		.out(chany_top_out[172]));

	mux_2level_tapbuf_size2 mux_top_track_346 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[174]}),
		.sram(mux_2level_tapbuf_size2_150_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_150_sram_inv[0:1]),
		.out(chany_top_out[173]));

	mux_2level_tapbuf_size2 mux_top_track_348 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[175]}),
		.sram(mux_2level_tapbuf_size2_151_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_151_sram_inv[0:1]),
		.out(chany_top_out[174]));

	mux_2level_tapbuf_size2 mux_top_track_350 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[176]}),
		.sram(mux_2level_tapbuf_size2_152_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_152_sram_inv[0:1]),
		.out(chany_top_out[175]));

	mux_2level_tapbuf_size2 mux_top_track_352 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[177]}),
		.sram(mux_2level_tapbuf_size2_153_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_153_sram_inv[0:1]),
		.out(chany_top_out[176]));

	mux_2level_tapbuf_size2 mux_top_track_354 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[178]}),
		.sram(mux_2level_tapbuf_size2_154_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_154_sram_inv[0:1]),
		.out(chany_top_out[177]));

	mux_2level_tapbuf_size2 mux_top_track_356 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[179]}),
		.sram(mux_2level_tapbuf_size2_155_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_155_sram_inv[0:1]),
		.out(chany_top_out[178]));

	mux_2level_tapbuf_size2 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[181]}),
		.sram(mux_2level_tapbuf_size2_156_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_156_sram_inv[0:1]),
		.out(chany_top_out[180]));

	mux_2level_tapbuf_size2 mux_top_track_362 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[182]}),
		.sram(mux_2level_tapbuf_size2_157_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_157_sram_inv[0:1]),
		.out(chany_top_out[181]));

	mux_2level_tapbuf_size2 mux_top_track_364 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[183]}),
		.sram(mux_2level_tapbuf_size2_158_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_158_sram_inv[0:1]),
		.out(chany_top_out[182]));

	mux_2level_tapbuf_size2 mux_top_track_366 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[184]}),
		.sram(mux_2level_tapbuf_size2_159_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_159_sram_inv[0:1]),
		.out(chany_top_out[183]));

	mux_2level_tapbuf_size2 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[185]}),
		.sram(mux_2level_tapbuf_size2_160_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_160_sram_inv[0:1]),
		.out(chany_top_out[184]));

	mux_2level_tapbuf_size2 mux_top_track_370 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[186]}),
		.sram(mux_2level_tapbuf_size2_161_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_161_sram_inv[0:1]),
		.out(chany_top_out[185]));

	mux_2level_tapbuf_size2 mux_top_track_372 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[187]}),
		.sram(mux_2level_tapbuf_size2_162_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_162_sram_inv[0:1]),
		.out(chany_top_out[186]));

	mux_2level_tapbuf_size2 mux_top_track_374 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[188]}),
		.sram(mux_2level_tapbuf_size2_163_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_163_sram_inv[0:1]),
		.out(chany_top_out[187]));

	mux_2level_tapbuf_size2 mux_top_track_378 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[190]}),
		.sram(mux_2level_tapbuf_size2_164_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_164_sram_inv[0:1]),
		.out(chany_top_out[189]));

	mux_2level_tapbuf_size2 mux_top_track_380 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[191]}),
		.sram(mux_2level_tapbuf_size2_165_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_165_sram_inv[0:1]),
		.out(chany_top_out[190]));

	mux_2level_tapbuf_size2 mux_top_track_382 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[192]}),
		.sram(mux_2level_tapbuf_size2_166_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_166_sram_inv[0:1]),
		.out(chany_top_out[191]));

	mux_2level_tapbuf_size2 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[193]}),
		.sram(mux_2level_tapbuf_size2_167_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_167_sram_inv[0:1]),
		.out(chany_top_out[192]));

	mux_2level_tapbuf_size2 mux_top_track_386 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[194]}),
		.sram(mux_2level_tapbuf_size2_168_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_168_sram_inv[0:1]),
		.out(chany_top_out[193]));

	mux_2level_tapbuf_size2 mux_top_track_388 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[195]}),
		.sram(mux_2level_tapbuf_size2_169_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_169_sram_inv[0:1]),
		.out(chany_top_out[194]));

	mux_2level_tapbuf_size2 mux_top_track_390 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[196]}),
		.sram(mux_2level_tapbuf_size2_170_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_170_sram_inv[0:1]),
		.out(chany_top_out[195]));

	mux_2level_tapbuf_size2 mux_top_track_392 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[197]}),
		.sram(mux_2level_tapbuf_size2_171_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_171_sram_inv[0:1]),
		.out(chany_top_out[196]));

	mux_2level_tapbuf_size2 mux_top_track_396 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[199]}),
		.sram(mux_2level_tapbuf_size2_172_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_172_sram_inv[0:1]),
		.out(chany_top_out[198]));

	mux_2level_tapbuf_size2 mux_top_track_398 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[200]}),
		.sram(mux_2level_tapbuf_size2_173_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_173_sram_inv[0:1]),
		.out(chany_top_out[199]));

	mux_2level_tapbuf_size2 mux_top_track_400 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[201]}),
		.sram(mux_2level_tapbuf_size2_174_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_174_sram_inv[0:1]),
		.out(chany_top_out[200]));

	mux_2level_tapbuf_size2 mux_top_track_402 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[202]}),
		.sram(mux_2level_tapbuf_size2_175_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_175_sram_inv[0:1]),
		.out(chany_top_out[201]));

	mux_2level_tapbuf_size2 mux_top_track_404 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[203]}),
		.sram(mux_2level_tapbuf_size2_176_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_176_sram_inv[0:1]),
		.out(chany_top_out[202]));

	mux_2level_tapbuf_size2 mux_top_track_406 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[204]}),
		.sram(mux_2level_tapbuf_size2_177_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_177_sram_inv[0:1]),
		.out(chany_top_out[203]));

	mux_2level_tapbuf_size2 mux_top_track_408 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[205]}),
		.sram(mux_2level_tapbuf_size2_178_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_178_sram_inv[0:1]),
		.out(chany_top_out[204]));

	mux_2level_tapbuf_size2 mux_top_track_410 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[206]}),
		.sram(mux_2level_tapbuf_size2_179_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_179_sram_inv[0:1]),
		.out(chany_top_out[205]));

	mux_2level_tapbuf_size2 mux_top_track_414 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[208]}),
		.sram(mux_2level_tapbuf_size2_180_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_180_sram_inv[0:1]),
		.out(chany_top_out[207]));

	mux_2level_tapbuf_size2 mux_top_track_416 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[209]}),
		.sram(mux_2level_tapbuf_size2_181_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_181_sram_inv[0:1]),
		.out(chany_top_out[208]));

	mux_2level_tapbuf_size2 mux_top_track_418 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[210]}),
		.sram(mux_2level_tapbuf_size2_182_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_182_sram_inv[0:1]),
		.out(chany_top_out[209]));

	mux_2level_tapbuf_size2 mux_top_track_420 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[211]}),
		.sram(mux_2level_tapbuf_size2_183_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_183_sram_inv[0:1]),
		.out(chany_top_out[210]));

	mux_2level_tapbuf_size2 mux_top_track_422 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[212]}),
		.sram(mux_2level_tapbuf_size2_184_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_184_sram_inv[0:1]),
		.out(chany_top_out[211]));

	mux_2level_tapbuf_size2 mux_top_track_424 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[213]}),
		.sram(mux_2level_tapbuf_size2_185_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_185_sram_inv[0:1]),
		.out(chany_top_out[212]));

	mux_2level_tapbuf_size2 mux_top_track_426 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[214]}),
		.sram(mux_2level_tapbuf_size2_186_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_186_sram_inv[0:1]),
		.out(chany_top_out[213]));

	mux_2level_tapbuf_size2 mux_top_track_428 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[215]}),
		.sram(mux_2level_tapbuf_size2_187_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_187_sram_inv[0:1]),
		.out(chany_top_out[214]));

	mux_2level_tapbuf_size2 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[217]}),
		.sram(mux_2level_tapbuf_size2_188_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_188_sram_inv[0:1]),
		.out(chany_top_out[216]));

	mux_2level_tapbuf_size2 mux_top_track_434 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[218]}),
		.sram(mux_2level_tapbuf_size2_189_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_189_sram_inv[0:1]),
		.out(chany_top_out[217]));

	mux_2level_tapbuf_size2 mux_top_track_436 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[219]}),
		.sram(mux_2level_tapbuf_size2_190_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_190_sram_inv[0:1]),
		.out(chany_top_out[218]));

	mux_2level_tapbuf_size2 mux_top_track_438 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[220]}),
		.sram(mux_2level_tapbuf_size2_191_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_191_sram_inv[0:1]),
		.out(chany_top_out[219]));

	mux_2level_tapbuf_size2 mux_top_track_440 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[221]}),
		.sram(mux_2level_tapbuf_size2_192_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_192_sram_inv[0:1]),
		.out(chany_top_out[220]));

	mux_2level_tapbuf_size2 mux_top_track_442 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[222]}),
		.sram(mux_2level_tapbuf_size2_193_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_193_sram_inv[0:1]),
		.out(chany_top_out[221]));

	mux_2level_tapbuf_size2 mux_top_track_444 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[223]}),
		.sram(mux_2level_tapbuf_size2_194_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_194_sram_inv[0:1]),
		.out(chany_top_out[222]));

	mux_2level_tapbuf_size2 mux_top_track_446 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[224]}),
		.sram(mux_2level_tapbuf_size2_195_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_195_sram_inv[0:1]),
		.out(chany_top_out[223]));

	mux_2level_tapbuf_size2 mux_top_track_450 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[226]}),
		.sram(mux_2level_tapbuf_size2_196_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_196_sram_inv[0:1]),
		.out(chany_top_out[225]));

	mux_2level_tapbuf_size2 mux_top_track_452 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[227]}),
		.sram(mux_2level_tapbuf_size2_197_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_197_sram_inv[0:1]),
		.out(chany_top_out[226]));

	mux_2level_tapbuf_size2 mux_top_track_454 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[228]}),
		.sram(mux_2level_tapbuf_size2_198_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_198_sram_inv[0:1]),
		.out(chany_top_out[227]));

	mux_2level_tapbuf_size2 mux_top_track_456 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[0]}),
		.sram(mux_2level_tapbuf_size2_199_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_199_sram_inv[0:1]),
		.out(chany_top_out[228]));

	mux_2level_tapbuf_size2 mux_right_track_8 (
		.in({chany_top_in[3], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_200_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_200_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size2 mux_right_track_10 (
		.in({chany_top_in[4], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_201_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_201_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size2 mux_right_track_12 (
		.in({chany_top_in[5], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_202_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_202_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size2 mux_right_track_14 (
		.in({chany_top_in[6], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_203_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_203_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size2 mux_right_track_18 (
		.in({chany_top_in[8], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_204_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_204_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size2 mux_right_track_20 (
		.in({chany_top_in[9], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_205_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_205_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size2 mux_right_track_22 (
		.in({chany_top_in[10], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_206_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_206_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size2 mux_right_track_24 (
		.in({chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_207_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_207_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size2 mux_right_track_26 (
		.in({chany_top_in[12], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_208_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_208_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size2 mux_right_track_28 (
		.in({chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_209_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_209_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size2 mux_right_track_30 (
		.in({chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_210_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_210_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size2 mux_right_track_32 (
		.in({chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_211_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_211_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size2 mux_right_track_36 (
		.in({chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_212_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_212_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size2 mux_right_track_38 (
		.in({chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_213_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_213_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size2 mux_right_track_40 (
		.in({chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_214_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_214_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size2 mux_right_track_42 (
		.in({chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_215_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_215_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size2 mux_right_track_44 (
		.in({chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_216_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_216_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size2 mux_right_track_46 (
		.in({chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_217_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_217_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size2 mux_right_track_48 (
		.in({chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_218_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_218_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size2 mux_right_track_50 (
		.in({chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_219_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_219_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size2 mux_right_track_54 (
		.in({chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_220_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_220_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size2 mux_right_track_56 (
		.in({chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_221_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_221_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size2 mux_right_track_58 (
		.in({chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_222_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_222_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size2 mux_right_track_60 (
		.in({chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_223_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_223_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size2 mux_right_track_62 (
		.in({chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_224_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_224_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size2 mux_right_track_64 (
		.in({chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_225_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_225_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size2 mux_right_track_66 (
		.in({chany_top_in[32], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_226_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_226_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size2 mux_right_track_68 (
		.in({chany_top_in[33], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_227_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_227_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size2 mux_right_track_72 (
		.in({chany_top_in[35], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_228_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_228_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size2 mux_right_track_74 (
		.in({chany_top_in[36], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_229_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_229_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size2 mux_right_track_76 (
		.in({chany_top_in[37], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_230_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_230_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size2 mux_right_track_78 (
		.in({chany_top_in[38], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_231_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_231_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size2 mux_right_track_80 (
		.in({chany_top_in[39], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_232_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_232_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size2 mux_right_track_82 (
		.in({chany_top_in[40], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_233_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_233_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size2 mux_right_track_84 (
		.in({chany_top_in[41], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_234_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_234_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size2 mux_right_track_86 (
		.in({chany_top_in[42], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_235_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_235_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size2 mux_right_track_90 (
		.in({chany_top_in[44], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_236_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_236_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size2 mux_right_track_92 (
		.in({chany_top_in[45], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_237_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_237_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size2 mux_right_track_94 (
		.in({chany_top_in[46], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_238_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_238_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size2 mux_right_track_96 (
		.in({chany_top_in[47], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_239_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_239_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size2 mux_right_track_98 (
		.in({chany_top_in[48], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_240_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_240_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size2 mux_right_track_100 (
		.in({chany_top_in[49], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_241_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_241_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size2 mux_right_track_102 (
		.in({chany_top_in[50], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_242_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_242_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size2 mux_right_track_104 (
		.in({chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_243_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_243_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size2 mux_right_track_108 (
		.in({chany_top_in[53], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_244_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_244_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size2 mux_right_track_110 (
		.in({chany_top_in[54], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_245_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_245_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size2 mux_right_track_112 (
		.in({chany_top_in[55], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_246_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_246_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size2 mux_right_track_114 (
		.in({chany_top_in[56], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_247_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_247_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size2 mux_right_track_116 (
		.in({chany_top_in[57], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_248_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_248_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size2 mux_right_track_118 (
		.in({chany_top_in[58], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_249_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_249_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_2level_tapbuf_size2 mux_right_track_120 (
		.in({chany_top_in[59], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_250_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_250_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size2 mux_right_track_122 (
		.in({chany_top_in[60], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_251_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_251_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size2 mux_right_track_126 (
		.in({chany_top_in[62], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_252_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_252_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size2 mux_right_track_128 (
		.in({chany_top_in[63], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_253_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_253_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size2 mux_right_track_130 (
		.in({chany_top_in[64], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_254_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_254_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size2 mux_right_track_132 (
		.in({chany_top_in[65], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_255_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_255_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size2 mux_right_track_134 (
		.in({chany_top_in[66], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_256_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_256_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size2 mux_right_track_136 (
		.in({chany_top_in[67], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_257_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_257_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size2 mux_right_track_138 (
		.in({chany_top_in[68], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_258_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_258_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size2 mux_right_track_140 (
		.in({chany_top_in[69], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_259_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_259_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size2 mux_right_track_144 (
		.in({chany_top_in[71], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_260_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_260_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size2 mux_right_track_146 (
		.in({chany_top_in[72], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_261_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_261_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size2 mux_right_track_148 (
		.in({chany_top_in[73], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_262_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_262_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size2 mux_right_track_150 (
		.in({chany_top_in[74], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_263_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_263_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size2 mux_right_track_152 (
		.in({chany_top_in[75], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_264_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_264_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size2 mux_right_track_154 (
		.in({chany_top_in[76], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_265_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_265_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size2 mux_right_track_156 (
		.in({chany_top_in[77], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_266_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_266_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size2 mux_right_track_158 (
		.in({chany_top_in[78], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_267_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_267_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_2level_tapbuf_size2 mux_right_track_162 (
		.in({chany_top_in[80], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_268_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_268_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size2 mux_right_track_164 (
		.in({chany_top_in[81], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_269_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_269_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size2 mux_right_track_166 (
		.in({chany_top_in[82], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_270_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_270_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size2 mux_right_track_168 (
		.in({chany_top_in[83], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_271_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_271_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size2 mux_right_track_170 (
		.in({chany_top_in[84], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_272_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_272_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size2 mux_right_track_172 (
		.in({chany_top_in[85], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_273_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_273_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size2 mux_right_track_174 (
		.in({chany_top_in[86], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_274_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_274_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size2 mux_right_track_176 (
		.in({chany_top_in[87], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_275_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_275_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size2 mux_right_track_180 (
		.in({chany_top_in[89], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_276_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_276_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size2 mux_right_track_182 (
		.in({chany_top_in[90], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_277_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_277_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size2 mux_right_track_184 (
		.in({chany_top_in[91], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_278_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_278_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size2 mux_right_track_186 (
		.in({chany_top_in[92], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_279_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_279_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size2 mux_right_track_188 (
		.in({chany_top_in[93], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_280_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_280_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size2 mux_right_track_190 (
		.in({chany_top_in[94], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_281_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_281_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size2 mux_right_track_192 (
		.in({chany_top_in[95], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_282_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_282_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size2 mux_right_track_194 (
		.in({chany_top_in[96], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_283_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_283_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size2 mux_right_track_198 (
		.in({chany_top_in[98], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_284_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_284_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_2level_tapbuf_size2 mux_right_track_200 (
		.in({chany_top_in[99], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_285_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_285_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size2 mux_right_track_202 (
		.in({chany_top_in[100], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_286_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_286_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size2 mux_right_track_204 (
		.in({chany_top_in[101], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_287_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_287_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size2 mux_right_track_206 (
		.in({chany_top_in[102], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_288_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_288_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_2level_tapbuf_size2 mux_right_track_208 (
		.in({chany_top_in[103], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_289_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_289_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size2 mux_right_track_210 (
		.in({chany_top_in[104], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_290_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_290_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size2 mux_right_track_212 (
		.in({chany_top_in[105], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_291_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_291_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size2 mux_right_track_216 (
		.in({chany_top_in[107], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_292_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_292_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size2 mux_right_track_218 (
		.in({chany_top_in[108], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_293_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_293_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_2level_tapbuf_size2 mux_right_track_220 (
		.in({chany_top_in[109], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_294_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_294_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size2 mux_right_track_222 (
		.in({chany_top_in[110], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_295_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_295_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_2level_tapbuf_size2 mux_right_track_224 (
		.in({chany_top_in[111], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_296_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_296_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size2 mux_right_track_226 (
		.in({chany_top_in[112], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_297_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_297_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size2 mux_right_track_228 (
		.in({chany_top_in[113], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_298_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_298_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size2 mux_right_track_230 (
		.in({chany_top_in[114], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_299_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_299_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_2level_tapbuf_size2 mux_right_track_234 (
		.in({chany_top_in[116], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_300_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_300_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size2 mux_right_track_236 (
		.in({chany_top_in[117], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_301_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_301_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_2level_tapbuf_size2 mux_right_track_238 (
		.in({chany_top_in[118], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_302_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_302_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_2level_tapbuf_size2 mux_right_track_240 (
		.in({chany_top_in[119], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_303_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_303_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size2 mux_right_track_242 (
		.in({chany_top_in[120], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_304_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_304_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size2 mux_right_track_244 (
		.in({chany_top_in[121], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_305_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_305_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size2 mux_right_track_246 (
		.in({chany_top_in[122], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_306_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_306_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_2level_tapbuf_size2 mux_right_track_248 (
		.in({chany_top_in[123], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_307_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_307_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size2 mux_right_track_252 (
		.in({chany_top_in[125], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_308_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_308_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size2 mux_right_track_254 (
		.in({chany_top_in[126], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_309_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_309_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_2level_tapbuf_size2 mux_right_track_256 (
		.in({chany_top_in[127], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_310_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_310_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size2 mux_right_track_258 (
		.in({chany_top_in[128], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_311_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_311_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_2level_tapbuf_size2 mux_right_track_260 (
		.in({chany_top_in[129], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_312_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_312_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size2 mux_right_track_262 (
		.in({chany_top_in[130], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_313_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_313_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_2level_tapbuf_size2 mux_right_track_264 (
		.in({chany_top_in[131], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_314_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_314_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size2 mux_right_track_266 (
		.in({chany_top_in[132], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_315_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_315_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size2 mux_right_track_270 (
		.in({chany_top_in[134], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_316_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_316_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_2level_tapbuf_size2 mux_right_track_272 (
		.in({chany_top_in[135], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_317_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_317_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size2 mux_right_track_274 (
		.in({chany_top_in[136], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_318_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_318_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size2 mux_right_track_276 (
		.in({chany_top_in[137], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_319_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_319_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_2level_tapbuf_size2 mux_right_track_278 (
		.in({chany_top_in[138], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_320_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_320_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_2level_tapbuf_size2 mux_right_track_280 (
		.in({chany_top_in[139], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_321_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_321_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size2 mux_right_track_282 (
		.in({chany_top_in[140], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_322_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_322_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size2 mux_right_track_284 (
		.in({chany_top_in[141], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_323_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_323_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size2 mux_right_track_288 (
		.in({chany_top_in[143], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_324_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_324_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size2 mux_right_track_290 (
		.in({chany_top_in[144], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_325_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_325_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size2 mux_right_track_292 (
		.in({chany_top_in[145], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_326_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_326_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size2 mux_right_track_294 (
		.in({chany_top_in[146], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_327_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_327_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_2level_tapbuf_size2 mux_right_track_296 (
		.in({chany_top_in[147], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_328_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_328_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size2 mux_right_track_298 (
		.in({chany_top_in[148], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_329_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_329_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_2level_tapbuf_size2 mux_right_track_300 (
		.in({chany_top_in[149], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_330_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_330_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_2level_tapbuf_size2 mux_right_track_302 (
		.in({chany_top_in[150], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_331_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_331_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_2level_tapbuf_size2 mux_right_track_306 (
		.in({chany_top_in[152], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_332_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_332_sram_inv[0:1]),
		.out(chanx_right_out[153]));

	mux_2level_tapbuf_size2 mux_right_track_308 (
		.in({chany_top_in[153], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_333_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_333_sram_inv[0:1]),
		.out(chanx_right_out[154]));

	mux_2level_tapbuf_size2 mux_right_track_310 (
		.in({chany_top_in[154], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_334_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_334_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_2level_tapbuf_size2 mux_right_track_312 (
		.in({chany_top_in[155], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_335_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_335_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_2level_tapbuf_size2 mux_right_track_314 (
		.in({chany_top_in[156], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_336_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_336_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_2level_tapbuf_size2 mux_right_track_316 (
		.in({chany_top_in[157], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_337_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_337_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_2level_tapbuf_size2 mux_right_track_318 (
		.in({chany_top_in[158], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_338_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_338_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_2level_tapbuf_size2 mux_right_track_320 (
		.in({chany_top_in[159], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_339_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_339_sram_inv[0:1]),
		.out(chanx_right_out[160]));

	mux_2level_tapbuf_size2 mux_right_track_324 (
		.in({chany_top_in[161], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_340_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_340_sram_inv[0:1]),
		.out(chanx_right_out[162]));

	mux_2level_tapbuf_size2 mux_right_track_326 (
		.in({chany_top_in[162], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_341_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_341_sram_inv[0:1]),
		.out(chanx_right_out[163]));

	mux_2level_tapbuf_size2 mux_right_track_328 (
		.in({chany_top_in[163], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_342_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_342_sram_inv[0:1]),
		.out(chanx_right_out[164]));

	mux_2level_tapbuf_size2 mux_right_track_330 (
		.in({chany_top_in[164], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_343_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_343_sram_inv[0:1]),
		.out(chanx_right_out[165]));

	mux_2level_tapbuf_size2 mux_right_track_332 (
		.in({chany_top_in[165], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_344_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_344_sram_inv[0:1]),
		.out(chanx_right_out[166]));

	mux_2level_tapbuf_size2 mux_right_track_334 (
		.in({chany_top_in[166], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_345_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_345_sram_inv[0:1]),
		.out(chanx_right_out[167]));

	mux_2level_tapbuf_size2 mux_right_track_336 (
		.in({chany_top_in[167], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_346_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_346_sram_inv[0:1]),
		.out(chanx_right_out[168]));

	mux_2level_tapbuf_size2 mux_right_track_338 (
		.in({chany_top_in[168], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_347_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_347_sram_inv[0:1]),
		.out(chanx_right_out[169]));

	mux_2level_tapbuf_size2 mux_right_track_342 (
		.in({chany_top_in[170], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_348_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_348_sram_inv[0:1]),
		.out(chanx_right_out[171]));

	mux_2level_tapbuf_size2 mux_right_track_344 (
		.in({chany_top_in[171], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_349_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_349_sram_inv[0:1]),
		.out(chanx_right_out[172]));

	mux_2level_tapbuf_size2 mux_right_track_346 (
		.in({chany_top_in[172], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_350_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_350_sram_inv[0:1]),
		.out(chanx_right_out[173]));

	mux_2level_tapbuf_size2 mux_right_track_348 (
		.in({chany_top_in[173], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_351_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_351_sram_inv[0:1]),
		.out(chanx_right_out[174]));

	mux_2level_tapbuf_size2 mux_right_track_350 (
		.in({chany_top_in[174], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_352_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_352_sram_inv[0:1]),
		.out(chanx_right_out[175]));

	mux_2level_tapbuf_size2 mux_right_track_352 (
		.in({chany_top_in[175], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_353_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_353_sram_inv[0:1]),
		.out(chanx_right_out[176]));

	mux_2level_tapbuf_size2 mux_right_track_354 (
		.in({chany_top_in[176], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_354_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_354_sram_inv[0:1]),
		.out(chanx_right_out[177]));

	mux_2level_tapbuf_size2 mux_right_track_356 (
		.in({chany_top_in[177], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_355_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_355_sram_inv[0:1]),
		.out(chanx_right_out[178]));

	mux_2level_tapbuf_size2 mux_right_track_360 (
		.in({chany_top_in[179], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_356_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_356_sram_inv[0:1]),
		.out(chanx_right_out[180]));

	mux_2level_tapbuf_size2 mux_right_track_362 (
		.in({chany_top_in[180], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_357_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_357_sram_inv[0:1]),
		.out(chanx_right_out[181]));

	mux_2level_tapbuf_size2 mux_right_track_364 (
		.in({chany_top_in[181], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_358_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_358_sram_inv[0:1]),
		.out(chanx_right_out[182]));

	mux_2level_tapbuf_size2 mux_right_track_366 (
		.in({chany_top_in[182], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_359_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_359_sram_inv[0:1]),
		.out(chanx_right_out[183]));

	mux_2level_tapbuf_size2 mux_right_track_368 (
		.in({chany_top_in[183], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_360_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_360_sram_inv[0:1]),
		.out(chanx_right_out[184]));

	mux_2level_tapbuf_size2 mux_right_track_370 (
		.in({chany_top_in[184], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_361_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_361_sram_inv[0:1]),
		.out(chanx_right_out[185]));

	mux_2level_tapbuf_size2 mux_right_track_372 (
		.in({chany_top_in[185], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_362_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_362_sram_inv[0:1]),
		.out(chanx_right_out[186]));

	mux_2level_tapbuf_size2 mux_right_track_374 (
		.in({chany_top_in[186], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_363_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_363_sram_inv[0:1]),
		.out(chanx_right_out[187]));

	mux_2level_tapbuf_size2 mux_right_track_378 (
		.in({chany_top_in[188], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_364_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_364_sram_inv[0:1]),
		.out(chanx_right_out[189]));

	mux_2level_tapbuf_size2 mux_right_track_380 (
		.in({chany_top_in[189], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_365_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_365_sram_inv[0:1]),
		.out(chanx_right_out[190]));

	mux_2level_tapbuf_size2 mux_right_track_382 (
		.in({chany_top_in[190], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_366_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_366_sram_inv[0:1]),
		.out(chanx_right_out[191]));

	mux_2level_tapbuf_size2 mux_right_track_384 (
		.in({chany_top_in[191], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_367_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_367_sram_inv[0:1]),
		.out(chanx_right_out[192]));

	mux_2level_tapbuf_size2 mux_right_track_386 (
		.in({chany_top_in[192], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_368_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_368_sram_inv[0:1]),
		.out(chanx_right_out[193]));

	mux_2level_tapbuf_size2 mux_right_track_388 (
		.in({chany_top_in[193], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_369_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_369_sram_inv[0:1]),
		.out(chanx_right_out[194]));

	mux_2level_tapbuf_size2 mux_right_track_390 (
		.in({chany_top_in[194], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_370_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_370_sram_inv[0:1]),
		.out(chanx_right_out[195]));

	mux_2level_tapbuf_size2 mux_right_track_392 (
		.in({chany_top_in[195], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_371_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_371_sram_inv[0:1]),
		.out(chanx_right_out[196]));

	mux_2level_tapbuf_size2 mux_right_track_396 (
		.in({chany_top_in[197], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_372_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_372_sram_inv[0:1]),
		.out(chanx_right_out[198]));

	mux_2level_tapbuf_size2 mux_right_track_398 (
		.in({chany_top_in[198], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_373_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_373_sram_inv[0:1]),
		.out(chanx_right_out[199]));

	mux_2level_tapbuf_size2 mux_right_track_400 (
		.in({chany_top_in[199], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_374_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_374_sram_inv[0:1]),
		.out(chanx_right_out[200]));

	mux_2level_tapbuf_size2 mux_right_track_402 (
		.in({chany_top_in[200], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_375_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_375_sram_inv[0:1]),
		.out(chanx_right_out[201]));

	mux_2level_tapbuf_size2 mux_right_track_404 (
		.in({chany_top_in[201], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_376_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_376_sram_inv[0:1]),
		.out(chanx_right_out[202]));

	mux_2level_tapbuf_size2 mux_right_track_406 (
		.in({chany_top_in[202], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_377_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_377_sram_inv[0:1]),
		.out(chanx_right_out[203]));

	mux_2level_tapbuf_size2 mux_right_track_408 (
		.in({chany_top_in[203], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_378_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_378_sram_inv[0:1]),
		.out(chanx_right_out[204]));

	mux_2level_tapbuf_size2 mux_right_track_410 (
		.in({chany_top_in[204], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_379_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_379_sram_inv[0:1]),
		.out(chanx_right_out[205]));

	mux_2level_tapbuf_size2 mux_right_track_414 (
		.in({chany_top_in[206], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_380_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_380_sram_inv[0:1]),
		.out(chanx_right_out[207]));

	mux_2level_tapbuf_size2 mux_right_track_416 (
		.in({chany_top_in[207], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_381_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_381_sram_inv[0:1]),
		.out(chanx_right_out[208]));

	mux_2level_tapbuf_size2 mux_right_track_418 (
		.in({chany_top_in[208], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_382_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_382_sram_inv[0:1]),
		.out(chanx_right_out[209]));

	mux_2level_tapbuf_size2 mux_right_track_420 (
		.in({chany_top_in[209], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_383_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_383_sram_inv[0:1]),
		.out(chanx_right_out[210]));

	mux_2level_tapbuf_size2 mux_right_track_422 (
		.in({chany_top_in[210], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_384_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_384_sram_inv[0:1]),
		.out(chanx_right_out[211]));

	mux_2level_tapbuf_size2 mux_right_track_424 (
		.in({chany_top_in[211], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_385_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_385_sram_inv[0:1]),
		.out(chanx_right_out[212]));

	mux_2level_tapbuf_size2 mux_right_track_426 (
		.in({chany_top_in[212], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_386_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_386_sram_inv[0:1]),
		.out(chanx_right_out[213]));

	mux_2level_tapbuf_size2 mux_right_track_428 (
		.in({chany_top_in[213], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_387_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_387_sram_inv[0:1]),
		.out(chanx_right_out[214]));

	mux_2level_tapbuf_size2 mux_right_track_432 (
		.in({chany_top_in[215], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_388_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_388_sram_inv[0:1]),
		.out(chanx_right_out[216]));

	mux_2level_tapbuf_size2 mux_right_track_434 (
		.in({chany_top_in[216], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_389_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_389_sram_inv[0:1]),
		.out(chanx_right_out[217]));

	mux_2level_tapbuf_size2 mux_right_track_436 (
		.in({chany_top_in[217], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_390_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_390_sram_inv[0:1]),
		.out(chanx_right_out[218]));

	mux_2level_tapbuf_size2 mux_right_track_438 (
		.in({chany_top_in[218], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_391_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_391_sram_inv[0:1]),
		.out(chanx_right_out[219]));

	mux_2level_tapbuf_size2 mux_right_track_440 (
		.in({chany_top_in[219], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_392_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_392_sram_inv[0:1]),
		.out(chanx_right_out[220]));

	mux_2level_tapbuf_size2 mux_right_track_442 (
		.in({chany_top_in[220], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_393_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_393_sram_inv[0:1]),
		.out(chanx_right_out[221]));

	mux_2level_tapbuf_size2 mux_right_track_444 (
		.in({chany_top_in[221], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_394_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_394_sram_inv[0:1]),
		.out(chanx_right_out[222]));

	mux_2level_tapbuf_size2 mux_right_track_446 (
		.in({chany_top_in[222], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_395_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_395_sram_inv[0:1]),
		.out(chanx_right_out[223]));

	mux_2level_tapbuf_size2 mux_right_track_450 (
		.in({chany_top_in[224], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_396_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_396_sram_inv[0:1]),
		.out(chanx_right_out[225]));

	mux_2level_tapbuf_size2 mux_right_track_452 (
		.in({chany_top_in[225], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_397_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_397_sram_inv[0:1]),
		.out(chanx_right_out[226]));

	mux_2level_tapbuf_size2 mux_right_track_454 (
		.in({chany_top_in[226], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_398_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_398_sram_inv[0:1]),
		.out(chanx_right_out[227]));

	mux_2level_tapbuf_size2 mux_right_track_456 (
		.in({chany_top_in[227], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_399_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_399_sram_inv[0:1]),
		.out(chanx_right_out[228]));

	mux_2level_tapbuf_size2_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_60_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_61_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_62_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_63_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_64_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_65_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_66_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_67_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_68_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_69_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_70_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_71_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_72_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_73_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_74_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_75_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_76_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_77_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_78_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_79_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_80_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_81_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_82_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_83_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_84_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_85_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_86_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_87_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_88_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_89_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_90_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_91_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_92_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_93_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_94_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_95_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_96_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_97_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_98_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_99_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_100_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_101_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_102_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_103_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_104_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_105_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_106_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_107_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_108_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_109_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_110_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_111_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_112_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_113_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_114_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_115_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_116_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_117_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_118_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_119_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_120_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_121_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_122_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_123_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_124_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_125_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_126_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_127_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_128_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_129_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_130_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_302 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_131_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_132_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_133_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_310 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_134_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_135_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_136_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_137_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_318 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_138_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_139_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_324 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_140_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_326 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_141_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_142_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_330 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_143_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_332 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_144_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_144_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_334 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_145_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_145_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_146_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_146_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_338 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_147_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_147_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_342 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_148_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_148_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_149_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_149_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_346 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_150_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_150_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_348 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_151_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_151_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_350 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_152_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_152_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_153_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_153_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_354 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_154_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_154_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_356 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_155_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_155_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_156_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_156_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_362 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_157_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_157_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_364 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_158_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_158_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_366 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_159_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_159_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_160_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_160_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_370 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_161_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_161_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_372 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_162_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_162_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_374 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_163_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_163_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_378 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_164_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_164_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_380 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_165_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_165_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_382 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_166_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_166_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_167_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_167_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_386 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_168_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_168_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_388 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_169_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_169_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_390 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_170_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_170_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_171_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_171_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_396 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_172_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_172_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_398 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_173_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_173_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_174_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_174_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_402 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_175_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_175_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_175_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_404 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_175_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_176_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_176_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_176_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_406 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_176_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_177_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_177_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_177_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_177_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_178_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_178_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_178_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_410 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_178_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_179_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_179_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_179_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_414 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_179_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_180_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_180_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_180_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_180_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_181_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_181_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_181_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_418 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_181_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_182_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_182_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_182_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_420 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_182_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_183_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_183_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_183_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_422 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_183_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_184_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_184_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_184_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_184_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_185_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_185_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_185_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_426 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_185_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_186_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_186_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_186_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_428 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_186_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_187_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_187_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_187_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_432 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_187_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_188_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_188_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_188_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_434 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_188_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_189_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_189_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_189_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_436 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_189_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_190_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_190_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_190_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_438 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_190_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_191_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_191_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_191_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_440 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_191_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_192_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_192_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_192_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_442 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_192_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_193_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_193_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_193_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_444 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_193_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_194_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_194_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_194_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_446 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_194_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_195_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_195_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_195_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_450 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_195_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_196_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_196_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_196_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_452 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_196_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_197_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_197_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_197_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_454 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_197_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_198_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_198_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_198_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_456 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_198_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_199_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_199_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_199_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_200_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_200_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_200_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_200_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_201_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_201_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_201_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_201_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_202_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_202_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_202_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_202_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_203_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_203_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_203_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_203_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_204_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_204_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_204_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_204_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_205_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_205_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_205_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_205_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_206_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_206_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_206_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_206_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_207_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_207_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_207_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_207_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_208_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_208_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_208_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_208_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_209_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_209_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_209_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_209_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_210_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_210_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_210_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_210_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_211_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_211_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_211_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_211_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_212_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_212_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_212_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_212_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_213_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_213_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_213_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_213_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_214_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_214_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_214_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_214_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_215_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_215_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_215_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_215_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_216_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_216_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_216_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_216_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_217_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_217_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_217_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_217_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_218_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_218_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_218_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_218_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_219_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_219_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_219_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_219_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_220_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_220_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_220_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_220_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_221_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_221_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_221_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_221_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_222_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_222_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_222_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_222_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_223_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_223_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_223_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_223_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_224_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_224_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_224_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_224_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_225_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_225_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_225_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_225_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_226_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_226_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_226_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_226_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_227_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_227_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_227_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_227_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_228_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_228_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_228_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_228_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_229_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_229_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_229_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_229_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_230_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_230_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_230_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_230_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_231_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_231_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_231_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_231_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_232_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_232_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_232_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_232_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_233_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_233_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_233_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_233_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_234_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_234_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_234_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_234_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_235_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_235_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_235_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_235_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_236_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_236_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_236_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_236_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_237_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_237_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_237_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_237_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_238_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_238_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_238_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_238_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_239_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_239_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_239_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_239_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_240_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_240_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_240_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_240_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_241_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_241_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_241_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_241_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_242_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_242_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_242_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_242_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_243_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_243_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_243_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_243_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_244_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_244_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_244_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_244_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_245_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_245_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_245_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_245_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_246_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_246_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_246_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_246_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_247_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_247_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_247_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_247_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_248_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_248_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_248_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_248_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_249_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_249_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_249_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_249_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_250_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_250_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_250_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_250_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_251_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_251_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_251_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_251_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_252_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_252_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_252_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_252_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_253_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_253_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_253_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_253_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_254_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_254_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_254_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_254_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_255_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_255_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_255_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_255_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_256_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_256_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_256_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_256_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_257_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_257_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_257_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_257_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_258_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_258_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_258_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_258_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_259_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_259_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_259_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_259_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_260_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_260_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_260_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_260_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_261_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_261_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_261_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_261_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_262_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_262_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_262_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_262_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_263_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_263_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_263_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_263_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_264_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_264_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_264_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_264_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_265_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_265_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_265_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_265_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_266_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_266_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_266_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_266_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_267_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_267_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_267_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_267_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_268_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_268_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_268_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_268_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_269_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_269_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_269_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_269_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_270_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_270_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_270_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_270_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_271_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_271_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_271_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_271_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_272_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_272_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_272_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_272_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_273_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_273_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_273_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_273_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_274_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_274_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_274_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_274_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_275_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_275_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_275_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_275_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_276_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_276_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_276_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_276_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_277_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_277_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_277_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_277_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_278_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_278_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_278_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_278_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_279_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_279_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_279_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_279_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_280_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_280_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_280_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_280_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_281_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_281_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_281_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_281_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_282_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_282_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_282_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_282_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_283_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_283_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_283_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_283_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_284_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_284_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_284_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_284_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_285_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_285_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_285_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_285_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_286_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_286_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_286_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_286_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_287_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_287_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_287_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_287_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_288_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_288_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_288_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_288_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_289_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_289_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_289_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_289_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_290_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_290_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_290_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_290_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_291_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_291_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_291_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_291_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_292_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_292_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_292_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_292_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_293_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_293_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_293_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_293_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_294_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_294_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_294_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_294_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_295_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_295_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_295_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_295_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_296_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_296_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_296_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_296_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_297_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_297_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_297_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_297_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_298_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_298_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_298_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_298_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_299_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_299_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_299_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_299_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_300_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_300_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_300_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_300_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_301_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_301_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_301_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_301_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_302_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_302_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_302_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_302_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_303_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_303_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_303_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_303_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_304_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_304_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_304_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_304_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_305_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_305_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_305_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_305_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_306_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_306_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_306_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_306_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_307_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_307_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_307_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_307_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_308_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_308_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_308_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_308_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_309_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_309_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_309_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_309_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_310_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_310_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_310_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_310_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_311_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_311_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_311_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_311_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_312_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_312_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_312_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_312_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_313_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_313_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_313_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_313_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_314_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_314_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_314_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_314_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_315_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_315_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_315_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_315_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_316_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_316_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_316_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_316_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_317_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_317_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_317_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_317_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_318_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_318_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_318_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_318_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_319_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_319_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_319_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_319_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_320_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_320_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_320_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_320_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_321_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_321_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_321_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_321_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_322_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_322_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_322_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_322_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_323_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_323_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_323_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_323_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_324_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_324_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_324_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_324_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_325_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_325_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_325_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_325_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_326_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_326_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_326_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_326_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_327_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_327_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_327_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_327_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_328_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_328_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_328_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_328_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_329_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_329_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_329_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_329_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_330_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_330_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_330_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_302 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_330_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_331_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_331_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_331_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_331_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_332_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_332_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_332_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_332_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_333_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_333_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_333_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_310 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_333_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_334_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_334_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_334_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_334_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_335_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_335_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_335_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_335_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_336_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_336_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_336_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_336_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_337_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_337_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_337_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_318 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_337_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_338_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_338_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_338_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_338_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_339_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_339_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_339_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_324 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_339_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_340_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_340_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_340_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_326 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_340_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_341_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_341_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_341_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_341_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_342_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_342_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_342_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_330 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_342_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_343_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_343_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_343_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_332 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_343_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_344_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_344_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_344_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_334 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_344_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_345_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_345_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_345_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_345_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_346_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_346_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_346_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_338 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_346_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_347_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_347_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_347_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_342 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_347_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_348_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_348_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_348_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_348_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_349_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_349_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_349_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_346 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_349_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_350_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_350_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_350_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_348 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_350_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_351_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_351_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_351_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_350 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_351_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_352_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_352_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_352_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_352_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_353_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_353_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_353_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_354 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_353_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_354_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_354_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_354_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_356 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_354_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_355_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_355_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_355_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_355_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_356_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_356_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_356_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_362 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_356_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_357_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_357_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_357_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_364 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_357_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_358_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_358_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_358_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_366 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_358_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_359_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_359_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_359_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_359_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_360_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_360_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_360_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_370 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_360_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_361_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_361_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_361_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_372 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_361_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_362_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_362_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_362_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_374 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_362_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_363_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_363_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_363_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_378 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_363_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_364_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_364_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_364_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_380 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_364_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_365_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_365_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_365_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_382 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_365_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_366_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_366_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_366_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_366_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_367_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_367_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_367_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_386 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_367_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_368_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_368_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_368_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_388 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_368_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_369_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_369_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_369_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_390 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_369_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_370_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_370_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_370_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_370_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_371_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_371_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_371_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_396 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_371_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_372_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_372_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_372_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_398 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_372_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_373_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_373_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_373_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_373_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_374_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_374_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_374_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_402 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_374_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_375_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_375_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_375_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_404 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_375_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_376_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_376_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_376_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_406 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_376_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_377_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_377_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_377_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_377_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_378_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_378_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_378_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_410 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_378_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_379_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_379_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_379_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_414 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_379_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_380_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_380_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_380_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_380_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_381_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_381_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_381_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_418 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_381_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_382_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_382_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_382_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_420 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_382_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_383_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_383_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_383_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_422 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_383_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_384_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_384_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_384_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_384_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_385_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_385_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_385_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_426 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_385_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_386_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_386_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_386_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_428 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_386_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_387_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_387_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_387_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_432 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_387_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_388_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_388_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_388_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_434 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_388_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_389_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_389_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_389_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_436 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_389_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_390_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_390_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_390_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_438 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_390_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_391_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_391_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_391_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_440 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_391_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_392_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_392_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_392_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_442 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_392_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_393_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_393_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_393_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_444 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_393_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_394_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_394_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_394_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_446 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_394_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_395_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_395_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_395_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_450 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_395_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_396_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_396_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_396_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_452 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_396_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_397_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_397_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_397_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_454 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_397_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_398_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_398_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_398_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_456 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_398_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_399_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_399_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__0_ -----

//----- Default net type -----
`default_nettype wire



