//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Oct 17 11:38:19 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__4_ -----
module sb_1__4_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:159] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:159] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_;
//----- INPUT PORTS -----
input [0:159] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:159] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:159] chany_top_out;
//----- OUTPUT PORTS -----
output [0:159] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:159] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:159] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size13_0_sram;
wire [0:7] mux_2level_tapbuf_size13_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_10_sram;
wire [0:7] mux_2level_tapbuf_size13_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_11_sram;
wire [0:7] mux_2level_tapbuf_size13_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_12_sram;
wire [0:7] mux_2level_tapbuf_size13_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_13_sram;
wire [0:7] mux_2level_tapbuf_size13_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_14_sram;
wire [0:7] mux_2level_tapbuf_size13_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_15_sram;
wire [0:7] mux_2level_tapbuf_size13_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_16_sram;
wire [0:7] mux_2level_tapbuf_size13_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_17_sram;
wire [0:7] mux_2level_tapbuf_size13_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_18_sram;
wire [0:7] mux_2level_tapbuf_size13_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_19_sram;
wire [0:7] mux_2level_tapbuf_size13_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_1_sram;
wire [0:7] mux_2level_tapbuf_size13_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_20_sram;
wire [0:7] mux_2level_tapbuf_size13_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_21_sram;
wire [0:7] mux_2level_tapbuf_size13_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_22_sram;
wire [0:7] mux_2level_tapbuf_size13_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_23_sram;
wire [0:7] mux_2level_tapbuf_size13_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_24_sram;
wire [0:7] mux_2level_tapbuf_size13_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_25_sram;
wire [0:7] mux_2level_tapbuf_size13_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_26_sram;
wire [0:7] mux_2level_tapbuf_size13_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_27_sram;
wire [0:7] mux_2level_tapbuf_size13_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_28_sram;
wire [0:7] mux_2level_tapbuf_size13_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_29_sram;
wire [0:7] mux_2level_tapbuf_size13_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_2_sram;
wire [0:7] mux_2level_tapbuf_size13_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_30_sram;
wire [0:7] mux_2level_tapbuf_size13_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_31_sram;
wire [0:7] mux_2level_tapbuf_size13_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_32_sram;
wire [0:7] mux_2level_tapbuf_size13_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_33_sram;
wire [0:7] mux_2level_tapbuf_size13_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_34_sram;
wire [0:7] mux_2level_tapbuf_size13_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_35_sram;
wire [0:7] mux_2level_tapbuf_size13_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_36_sram;
wire [0:7] mux_2level_tapbuf_size13_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_37_sram;
wire [0:7] mux_2level_tapbuf_size13_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_38_sram;
wire [0:7] mux_2level_tapbuf_size13_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_39_sram;
wire [0:7] mux_2level_tapbuf_size13_39_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_3_sram;
wire [0:7] mux_2level_tapbuf_size13_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_40_sram;
wire [0:7] mux_2level_tapbuf_size13_40_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_41_sram;
wire [0:7] mux_2level_tapbuf_size13_41_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_42_sram;
wire [0:7] mux_2level_tapbuf_size13_42_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_43_sram;
wire [0:7] mux_2level_tapbuf_size13_43_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_44_sram;
wire [0:7] mux_2level_tapbuf_size13_44_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_45_sram;
wire [0:7] mux_2level_tapbuf_size13_45_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_46_sram;
wire [0:7] mux_2level_tapbuf_size13_46_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_47_sram;
wire [0:7] mux_2level_tapbuf_size13_47_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_48_sram;
wire [0:7] mux_2level_tapbuf_size13_48_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_49_sram;
wire [0:7] mux_2level_tapbuf_size13_49_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_4_sram;
wire [0:7] mux_2level_tapbuf_size13_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_50_sram;
wire [0:7] mux_2level_tapbuf_size13_50_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_51_sram;
wire [0:7] mux_2level_tapbuf_size13_51_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_52_sram;
wire [0:7] mux_2level_tapbuf_size13_52_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_53_sram;
wire [0:7] mux_2level_tapbuf_size13_53_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_54_sram;
wire [0:7] mux_2level_tapbuf_size13_54_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_55_sram;
wire [0:7] mux_2level_tapbuf_size13_55_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_56_sram;
wire [0:7] mux_2level_tapbuf_size13_56_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_57_sram;
wire [0:7] mux_2level_tapbuf_size13_57_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_58_sram;
wire [0:7] mux_2level_tapbuf_size13_58_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_59_sram;
wire [0:7] mux_2level_tapbuf_size13_59_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_5_sram;
wire [0:7] mux_2level_tapbuf_size13_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_60_sram;
wire [0:7] mux_2level_tapbuf_size13_60_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_61_sram;
wire [0:7] mux_2level_tapbuf_size13_61_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_62_sram;
wire [0:7] mux_2level_tapbuf_size13_62_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_63_sram;
wire [0:7] mux_2level_tapbuf_size13_63_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_64_sram;
wire [0:7] mux_2level_tapbuf_size13_64_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_65_sram;
wire [0:7] mux_2level_tapbuf_size13_65_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_66_sram;
wire [0:7] mux_2level_tapbuf_size13_66_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_67_sram;
wire [0:7] mux_2level_tapbuf_size13_67_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_68_sram;
wire [0:7] mux_2level_tapbuf_size13_68_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_69_sram;
wire [0:7] mux_2level_tapbuf_size13_69_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_6_sram;
wire [0:7] mux_2level_tapbuf_size13_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_70_sram;
wire [0:7] mux_2level_tapbuf_size13_70_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_71_sram;
wire [0:7] mux_2level_tapbuf_size13_71_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_72_sram;
wire [0:7] mux_2level_tapbuf_size13_72_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_73_sram;
wire [0:7] mux_2level_tapbuf_size13_73_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_74_sram;
wire [0:7] mux_2level_tapbuf_size13_74_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_75_sram;
wire [0:7] mux_2level_tapbuf_size13_75_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_76_sram;
wire [0:7] mux_2level_tapbuf_size13_76_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_77_sram;
wire [0:7] mux_2level_tapbuf_size13_77_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_78_sram;
wire [0:7] mux_2level_tapbuf_size13_78_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_79_sram;
wire [0:7] mux_2level_tapbuf_size13_79_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_7_sram;
wire [0:7] mux_2level_tapbuf_size13_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_8_sram;
wire [0:7] mux_2level_tapbuf_size13_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_9_sram;
wire [0:7] mux_2level_tapbuf_size13_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_9_ccff_tail;
wire [0:11] mux_2level_tapbuf_size25_0_sram;
wire [0:11] mux_2level_tapbuf_size25_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size25_mem_0_ccff_tail;
wire [0:11] mux_2level_tapbuf_size26_0_sram;
wire [0:11] mux_2level_tapbuf_size26_0_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_10_sram;
wire [0:11] mux_2level_tapbuf_size26_10_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_11_sram;
wire [0:11] mux_2level_tapbuf_size26_11_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_12_sram;
wire [0:11] mux_2level_tapbuf_size26_12_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_13_sram;
wire [0:11] mux_2level_tapbuf_size26_13_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_14_sram;
wire [0:11] mux_2level_tapbuf_size26_14_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_15_sram;
wire [0:11] mux_2level_tapbuf_size26_15_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_16_sram;
wire [0:11] mux_2level_tapbuf_size26_16_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_17_sram;
wire [0:11] mux_2level_tapbuf_size26_17_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_18_sram;
wire [0:11] mux_2level_tapbuf_size26_18_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_19_sram;
wire [0:11] mux_2level_tapbuf_size26_19_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_1_sram;
wire [0:11] mux_2level_tapbuf_size26_1_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_20_sram;
wire [0:11] mux_2level_tapbuf_size26_20_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_21_sram;
wire [0:11] mux_2level_tapbuf_size26_21_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_22_sram;
wire [0:11] mux_2level_tapbuf_size26_22_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_23_sram;
wire [0:11] mux_2level_tapbuf_size26_23_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_24_sram;
wire [0:11] mux_2level_tapbuf_size26_24_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_25_sram;
wire [0:11] mux_2level_tapbuf_size26_25_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_26_sram;
wire [0:11] mux_2level_tapbuf_size26_26_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_27_sram;
wire [0:11] mux_2level_tapbuf_size26_27_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_28_sram;
wire [0:11] mux_2level_tapbuf_size26_28_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_29_sram;
wire [0:11] mux_2level_tapbuf_size26_29_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_2_sram;
wire [0:11] mux_2level_tapbuf_size26_2_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_30_sram;
wire [0:11] mux_2level_tapbuf_size26_30_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_3_sram;
wire [0:11] mux_2level_tapbuf_size26_3_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_4_sram;
wire [0:11] mux_2level_tapbuf_size26_4_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_5_sram;
wire [0:11] mux_2level_tapbuf_size26_5_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_6_sram;
wire [0:11] mux_2level_tapbuf_size26_6_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_7_sram;
wire [0:11] mux_2level_tapbuf_size26_7_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_8_sram;
wire [0:11] mux_2level_tapbuf_size26_8_sram_inv;
wire [0:11] mux_2level_tapbuf_size26_9_sram;
wire [0:11] mux_2level_tapbuf_size26_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size26_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size26_mem_9_ccff_tail;
wire [0:11] mux_2level_tapbuf_size27_0_sram;
wire [0:11] mux_2level_tapbuf_size27_0_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_1_sram;
wire [0:11] mux_2level_tapbuf_size27_1_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_2_sram;
wire [0:11] mux_2level_tapbuf_size27_2_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_3_sram;
wire [0:11] mux_2level_tapbuf_size27_3_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_4_sram;
wire [0:11] mux_2level_tapbuf_size27_4_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_5_sram;
wire [0:11] mux_2level_tapbuf_size27_5_sram_inv;
wire [0:11] mux_2level_tapbuf_size27_6_sram;
wire [0:11] mux_2level_tapbuf_size27_6_sram_inv;
wire [0:0] mux_2level_tapbuf_size27_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size27_mem_6_ccff_tail;
wire [0:11] mux_2level_tapbuf_size29_0_sram;
wire [0:11] mux_2level_tapbuf_size29_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size29_mem_0_ccff_tail;
wire [0:13] mux_2level_tapbuf_size42_0_sram;
wire [0:13] mux_2level_tapbuf_size42_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size42_mem_0_ccff_tail;
wire [0:13] mux_2level_tapbuf_size43_0_sram;
wire [0:13] mux_2level_tapbuf_size43_0_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_10_sram;
wire [0:13] mux_2level_tapbuf_size43_10_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_11_sram;
wire [0:13] mux_2level_tapbuf_size43_11_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_12_sram;
wire [0:13] mux_2level_tapbuf_size43_12_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_13_sram;
wire [0:13] mux_2level_tapbuf_size43_13_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_14_sram;
wire [0:13] mux_2level_tapbuf_size43_14_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_15_sram;
wire [0:13] mux_2level_tapbuf_size43_15_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_16_sram;
wire [0:13] mux_2level_tapbuf_size43_16_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_17_sram;
wire [0:13] mux_2level_tapbuf_size43_17_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_18_sram;
wire [0:13] mux_2level_tapbuf_size43_18_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_19_sram;
wire [0:13] mux_2level_tapbuf_size43_19_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_1_sram;
wire [0:13] mux_2level_tapbuf_size43_1_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_20_sram;
wire [0:13] mux_2level_tapbuf_size43_20_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_21_sram;
wire [0:13] mux_2level_tapbuf_size43_21_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_22_sram;
wire [0:13] mux_2level_tapbuf_size43_22_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_2_sram;
wire [0:13] mux_2level_tapbuf_size43_2_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_3_sram;
wire [0:13] mux_2level_tapbuf_size43_3_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_4_sram;
wire [0:13] mux_2level_tapbuf_size43_4_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_5_sram;
wire [0:13] mux_2level_tapbuf_size43_5_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_6_sram;
wire [0:13] mux_2level_tapbuf_size43_6_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_7_sram;
wire [0:13] mux_2level_tapbuf_size43_7_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_8_sram;
wire [0:13] mux_2level_tapbuf_size43_8_sram_inv;
wire [0:13] mux_2level_tapbuf_size43_9_sram;
wire [0:13] mux_2level_tapbuf_size43_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size43_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size43_mem_9_ccff_tail;
wire [0:13] mux_2level_tapbuf_size44_0_sram;
wire [0:13] mux_2level_tapbuf_size44_0_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_10_sram;
wire [0:13] mux_2level_tapbuf_size44_10_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_11_sram;
wire [0:13] mux_2level_tapbuf_size44_11_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_12_sram;
wire [0:13] mux_2level_tapbuf_size44_12_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_13_sram;
wire [0:13] mux_2level_tapbuf_size44_13_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_14_sram;
wire [0:13] mux_2level_tapbuf_size44_14_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_1_sram;
wire [0:13] mux_2level_tapbuf_size44_1_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_2_sram;
wire [0:13] mux_2level_tapbuf_size44_2_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_3_sram;
wire [0:13] mux_2level_tapbuf_size44_3_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_4_sram;
wire [0:13] mux_2level_tapbuf_size44_4_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_5_sram;
wire [0:13] mux_2level_tapbuf_size44_5_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_6_sram;
wire [0:13] mux_2level_tapbuf_size44_6_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_7_sram;
wire [0:13] mux_2level_tapbuf_size44_7_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_8_sram;
wire [0:13] mux_2level_tapbuf_size44_8_sram_inv;
wire [0:13] mux_2level_tapbuf_size44_9_sram;
wire [0:13] mux_2level_tapbuf_size44_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size44_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size44_mem_9_ccff_tail;
wire [0:13] mux_2level_tapbuf_size46_0_sram;
wire [0:13] mux_2level_tapbuf_size46_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size46_mem_0_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[64] = chany_top_in[64];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[68] = chany_top_in[68];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[72] = chany_top_in[72];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[76] = chany_top_in[76];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[80] = chany_top_in[80];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[84] = chany_top_in[84];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[88] = chany_top_in[88];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[92] = chany_top_in[92];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[96] = chany_top_in[96];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[98];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[100] = chany_top_in[100];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[102];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[104] = chany_top_in[104];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[106];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[108] = chany_top_in[108];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[110];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[112] = chany_top_in[112];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[114];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[116] = chany_top_in[116];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[118];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[120] = chany_top_in[120];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[122];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[124] = chany_top_in[124];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[126];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[128] = chany_top_in[128];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[130];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[132] = chany_top_in[132];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[134];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[136] = chany_top_in[136];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[138];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[140] = chany_top_in[140];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[142];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[144] = chany_top_in[144];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[146];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[148] = chany_top_in[148];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[150];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[152] = chany_top_in[152];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[154];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[156] = chany_top_in[156];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[158];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[159];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[0] = chanx_right_in[0];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[2];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[3];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[4] = chanx_right_in[4];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[6];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[7];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[8] = chanx_right_in[8];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[10];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[11];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[12] = chanx_right_in[12];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[14];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[15];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[16] = chanx_right_in[16];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[18];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[19];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[20] = chanx_right_in[20];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[22];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[23];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[24] = chanx_right_in[24];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[26];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[27];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[28] = chanx_right_in[28];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[30];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[31];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[64] = chanx_right_in[64];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[66] = chanx_right_in[66];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[67] = chanx_right_in[67];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[68] = chanx_right_in[68];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[70] = chanx_right_in[70];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[71] = chanx_right_in[71];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[72] = chanx_right_in[72];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[74] = chanx_right_in[74];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[75] = chanx_right_in[75];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[76] = chanx_right_in[76];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[78] = chanx_right_in[78];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[79];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[80] = chanx_right_in[80];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[82];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[83];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[84] = chanx_right_in[84];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[86];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[87];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[88] = chanx_right_in[88];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[90] = chanx_right_in[90];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[91];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[92] = chanx_right_in[92];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[94] = chanx_right_in[94];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[95];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[96] = chanx_right_in[96];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[98] = chanx_right_in[98];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[99];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[100] = chanx_right_in[100];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[102] = chanx_right_in[102];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[103] = chanx_right_in[103];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[104] = chanx_right_in[104];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[106] = chanx_right_in[106];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[107] = chanx_right_in[107];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[108] = chanx_right_in[108];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[110] = chanx_right_in[110];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[111] = chanx_right_in[111];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[112] = chanx_right_in[112];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[114] = chanx_right_in[114];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[115] = chanx_right_in[115];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[116] = chanx_right_in[116];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[118] = chanx_right_in[118];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[119] = chanx_right_in[119];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[120] = chanx_right_in[120];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[122] = chanx_right_in[122];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[123] = chanx_right_in[123];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[124] = chanx_right_in[124];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[126] = chanx_right_in[126];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[127] = chanx_right_in[127];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[128] = chanx_right_in[128];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[130] = chanx_right_in[130];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[131] = chanx_right_in[131];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[132] = chanx_right_in[132];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[134] = chanx_right_in[134];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[135] = chanx_right_in[135];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[136] = chanx_right_in[136];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[138] = chanx_right_in[138];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[139] = chanx_right_in[139];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[140] = chanx_right_in[140];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[142] = chanx_right_in[142];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[143] = chanx_right_in[143];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[144] = chanx_right_in[144];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[146] = chanx_right_in[146];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[147] = chanx_right_in[147];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[148] = chanx_right_in[148];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[150] = chanx_right_in[150];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[151] = chanx_right_in[151];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[152] = chanx_right_in[152];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[154] = chanx_right_in[154];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[155] = chanx_right_in[155];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[156] = chanx_right_in[156];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[158] = chanx_right_in[158];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[159] = chanx_right_in[159];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[2];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[6];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[10];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[14];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[18];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[22];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[26];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[30];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[34];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[38];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[42];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[46];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[50];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[54];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[58];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[62];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[64];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[66];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[67];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[68];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[70];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[71];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chany_bottom_in[72];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[74];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[75];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chany_bottom_in[76];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[78];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[79];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chany_bottom_in[80];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[82];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[83];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chany_bottom_in[84];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[86];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[87];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chany_bottom_in[88];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[90];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[91];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chany_bottom_in[92];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[94];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[95];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[96] = chany_bottom_in[96];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[98];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[99];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[100] = chany_bottom_in[100];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[102];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[103];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[104] = chany_bottom_in[104];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[106];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[107];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[108] = chany_bottom_in[108];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[110];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[111];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[112] = chany_bottom_in[112];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[114];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[115];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chany_bottom_in[116];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[118];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[119];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[120] = chany_bottom_in[120];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[122];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[123];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[124] = chany_bottom_in[124];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[126];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[127];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[128] = chany_bottom_in[128];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[130];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[131];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chany_bottom_in[132];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[134];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[135];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[136] = chany_bottom_in[136];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[138];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[139];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[140] = chany_bottom_in[140];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[142];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[143];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[144] = chany_bottom_in[144];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[146];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[147];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[148] = chany_bottom_in[148];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[150];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[151];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chany_bottom_in[152];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[154];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[155];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[156] = chany_bottom_in[156];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[158];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[159];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[0] = chanx_left_in[0];
// ----- Local connection due to Wire 631 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[2];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[3];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[4] = chanx_left_in[4];
// ----- Local connection due to Wire 635 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[6];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[7];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[8] = chanx_left_in[8];
// ----- Local connection due to Wire 639 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[10];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[11];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[12] = chanx_left_in[12];
// ----- Local connection due to Wire 643 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[14];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[15];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[16] = chanx_left_in[16];
// ----- Local connection due to Wire 647 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[18];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[19];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[20] = chanx_left_in[20];
// ----- Local connection due to Wire 651 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[22];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[23];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[24] = chanx_left_in[24];
// ----- Local connection due to Wire 655 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[26];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[27];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[28] = chanx_left_in[28];
// ----- Local connection due to Wire 659 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[30];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[31];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 663 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[34];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 667 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[38];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 671 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[42];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 675 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[46];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 679 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[50];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 683 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[54];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 687 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[58];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 691 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[62];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[64] = chanx_left_in[64];
// ----- Local connection due to Wire 695 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[66];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[67];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[68] = chanx_left_in[68];
// ----- Local connection due to Wire 699 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[70];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[71];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[72] = chanx_left_in[72];
// ----- Local connection due to Wire 703 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[74];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[75];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[76] = chanx_left_in[76];
// ----- Local connection due to Wire 707 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[78];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[79];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[80] = chanx_left_in[80];
// ----- Local connection due to Wire 711 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[82];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[83];
// ----- Local connection due to Wire 713 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[84] = chanx_left_in[84];
// ----- Local connection due to Wire 715 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[86];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[87];
// ----- Local connection due to Wire 717 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[88] = chanx_left_in[88];
// ----- Local connection due to Wire 719 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[90];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[91];
// ----- Local connection due to Wire 721 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[92] = chanx_left_in[92];
// ----- Local connection due to Wire 723 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[94];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[95];
// ----- Local connection due to Wire 725 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[96] = chanx_left_in[96];
// ----- Local connection due to Wire 727 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[98];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[99];
// ----- Local connection due to Wire 729 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[100] = chanx_left_in[100];
// ----- Local connection due to Wire 731 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[102];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[103];
// ----- Local connection due to Wire 733 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[104] = chanx_left_in[104];
// ----- Local connection due to Wire 735 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[106];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[107];
// ----- Local connection due to Wire 737 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[108] = chanx_left_in[108];
// ----- Local connection due to Wire 739 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[110];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[111];
// ----- Local connection due to Wire 741 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[112] = chanx_left_in[112];
// ----- Local connection due to Wire 743 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[114];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[115];
// ----- Local connection due to Wire 745 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[116] = chanx_left_in[116];
// ----- Local connection due to Wire 747 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[118];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[119];
// ----- Local connection due to Wire 749 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[120] = chanx_left_in[120];
// ----- Local connection due to Wire 751 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[122];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[123];
// ----- Local connection due to Wire 753 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[124] = chanx_left_in[124];
// ----- Local connection due to Wire 755 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[126];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[127];
// ----- Local connection due to Wire 757 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[128] = chanx_left_in[128];
// ----- Local connection due to Wire 759 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[130];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[131];
// ----- Local connection due to Wire 761 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[132] = chanx_left_in[132];
// ----- Local connection due to Wire 763 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[134];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[135];
// ----- Local connection due to Wire 765 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[136] = chanx_left_in[136];
// ----- Local connection due to Wire 767 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[138];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[139];
// ----- Local connection due to Wire 769 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[140] = chanx_left_in[140];
// ----- Local connection due to Wire 771 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[142];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[143];
// ----- Local connection due to Wire 773 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[144] = chanx_left_in[144];
// ----- Local connection due to Wire 775 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[146];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[147];
// ----- Local connection due to Wire 777 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[148] = chanx_left_in[148];
// ----- Local connection due to Wire 779 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[150];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[151];
// ----- Local connection due to Wire 781 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[152] = chanx_left_in[152];
// ----- Local connection due to Wire 783 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[154];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[155];
// ----- Local connection due to Wire 785 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[156] = chanx_left_in[156];
// ----- Local connection due to Wire 787 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[158];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[159];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size13 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[2], chanx_right_in[5], chanx_right_in[55], chanx_right_in[108], chany_bottom_in[1], chanx_left_in[0:1], chanx_left_in[54], chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size13_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_0_sram_inv[0:7]),
		.out(chany_top_out[1]));

	mux_2level_tapbuf_size13 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[3], chanx_right_in[9], chanx_right_in[56], chanx_right_in[110], chany_bottom_in[5], chanx_left_in[52], chanx_left_in[106], chanx_left_in[157], chanx_left_in[159]}),
		.sram(mux_2level_tapbuf_size13_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_1_sram_inv[0:7]),
		.out(chany_top_out[5]));

	mux_2level_tapbuf_size13 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[4], chanx_right_in[13], chanx_right_in[58], chanx_right_in[111], chany_bottom_in[9], chanx_left_in[51], chanx_left_in[104], chanx_left_in[153], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size13_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_2_sram_inv[0:7]),
		.out(chany_top_out[9]));

	mux_2level_tapbuf_size13 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[6], chanx_right_in[17], chanx_right_in[59], chanx_right_in[112], chany_bottom_in[13], chanx_left_in[50], chanx_left_in[103], chanx_left_in[149], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size13_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_3_sram_inv[0:7]),
		.out(chany_top_out[13]));

	mux_2level_tapbuf_size13 mux_top_track_34 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[7], chanx_right_in[21], chanx_right_in[60], chanx_right_in[114], chany_bottom_in[17], chanx_left_in[48], chanx_left_in[102], chanx_left_in[145], chanx_left_in[155]}),
		.sram(mux_2level_tapbuf_size13_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_4_sram_inv[0:7]),
		.out(chany_top_out[17]));

	mux_2level_tapbuf_size13 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[8], chanx_right_in[25], chanx_right_in[62], chanx_right_in[115], chany_bottom_in[21], chanx_left_in[47], chanx_left_in[100], chanx_left_in[141], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size13_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_5_sram_inv[0:7]),
		.out(chany_top_out[21]));

	mux_2level_tapbuf_size13 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[10], chanx_right_in[29], chanx_right_in[63], chanx_right_in[116], chany_bottom_in[25], chanx_left_in[46], chanx_left_in[99], chanx_left_in[137], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size13_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_6_sram_inv[0:7]),
		.out(chany_top_out[25]));

	mux_2level_tapbuf_size13 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[11], chanx_right_in[33], chanx_right_in[64], chanx_right_in[118], chany_bottom_in[29], chanx_left_in[44], chanx_left_in[98], chanx_left_in[133], chanx_left_in[151]}),
		.sram(mux_2level_tapbuf_size13_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_7_sram_inv[0:7]),
		.out(chany_top_out[29]));

	mux_2level_tapbuf_size13 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[12], chanx_right_in[37], chanx_right_in[66], chanx_right_in[119], chany_bottom_in[33], chanx_left_in[43], chanx_left_in[96], chanx_left_in[129], chanx_left_in[150]}),
		.sram(mux_2level_tapbuf_size13_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_8_sram_inv[0:7]),
		.out(chany_top_out[33]));

	mux_2level_tapbuf_size13 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[14], chanx_right_in[41], chanx_right_in[67], chanx_right_in[120], chany_bottom_in[37], chanx_left_in[42], chanx_left_in[95], chanx_left_in[125], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size13_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_9_sram_inv[0:7]),
		.out(chany_top_out[37]));

	mux_2level_tapbuf_size13 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[15], chanx_right_in[45], chanx_right_in[68], chanx_right_in[122], chany_bottom_in[41], chanx_left_in[40], chanx_left_in[94], chanx_left_in[121], chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size13_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_10_sram_inv[0:7]),
		.out(chany_top_out[41]));

	mux_2level_tapbuf_size13 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[16], chanx_right_in[49], chanx_right_in[70], chanx_right_in[123], chany_bottom_in[45], chanx_left_in[39], chanx_left_in[92], chanx_left_in[117], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size13_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_11_sram_inv[0:7]),
		.out(chany_top_out[45]));

	mux_2level_tapbuf_size13 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[18], chanx_right_in[53], chanx_right_in[71], chanx_right_in[124], chany_bottom_in[49], chanx_left_in[38], chanx_left_in[91], chanx_left_in[113], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size13_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_12_sram_inv[0:7]),
		.out(chany_top_out[49]));

	mux_2level_tapbuf_size13 mux_top_track_106 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[19], chanx_right_in[57], chanx_right_in[72], chanx_right_in[126], chany_bottom_in[53], chanx_left_in[36], chanx_left_in[90], chanx_left_in[109], chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size13_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_13_sram_inv[0:7]),
		.out(chany_top_out[53]));

	mux_2level_tapbuf_size13 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[20], chanx_right_in[61], chanx_right_in[74], chanx_right_in[127], chany_bottom_in[57], chanx_left_in[35], chanx_left_in[88], chanx_left_in[105], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size13_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_14_sram_inv[0:7]),
		.out(chany_top_out[57]));

	mux_2level_tapbuf_size13 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[22], chanx_right_in[65], chanx_right_in[75], chanx_right_in[128], chany_bottom_in[61], chanx_left_in[34], chanx_left_in[87], chanx_left_in[101], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size13_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_15_sram_inv[0:7]),
		.out(chany_top_out[61]));

	mux_2level_tapbuf_size13 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[23], chanx_right_in[69], chanx_right_in[76], chanx_right_in[130], chany_bottom_in[65], chanx_left_in[32], chanx_left_in[86], chanx_left_in[97], chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size13_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_16_sram_inv[0:7]),
		.out(chany_top_out[65]));

	mux_2level_tapbuf_size13 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[24], chanx_right_in[73], chanx_right_in[78], chanx_right_in[131], chany_bottom_in[69], chanx_left_in[31], chanx_left_in[84], chanx_left_in[93], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size13_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_17_sram_inv[0:7]),
		.out(chany_top_out[69]));

	mux_2level_tapbuf_size13 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[26], chanx_right_in[77], chanx_right_in[79], chanx_right_in[132], chany_bottom_in[73], chanx_left_in[30], chanx_left_in[83], chanx_left_in[89], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size13_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_18_sram_inv[0:7]),
		.out(chany_top_out[73]));

	mux_2level_tapbuf_size13 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[27], chanx_right_in[80:81], chanx_right_in[134], chany_bottom_in[77], chanx_left_in[28], chanx_left_in[82], chanx_left_in[85], chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size13_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_19_sram_inv[0:7]),
		.out(chany_top_out[77]));

	mux_2level_tapbuf_size13 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[28], chanx_right_in[82], chanx_right_in[85], chanx_right_in[135], chany_bottom_in[81], chanx_left_in[27], chanx_left_in[80:81], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size13_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_20_sram_inv[0:7]),
		.out(chany_top_out[81]));

	mux_2level_tapbuf_size13 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[30], chanx_right_in[83], chanx_right_in[89], chanx_right_in[136], chany_bottom_in[85], chanx_left_in[26], chanx_left_in[77], chanx_left_in[79], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size13_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_21_sram_inv[0:7]),
		.out(chany_top_out[85]));

	mux_2level_tapbuf_size13 mux_top_track_178 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[31], chanx_right_in[84], chanx_right_in[93], chanx_right_in[138], chany_bottom_in[89], chanx_left_in[24], chanx_left_in[73], chanx_left_in[78], chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size13_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_22_sram_inv[0:7]),
		.out(chany_top_out[89]));

	mux_2level_tapbuf_size13 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[32], chanx_right_in[86], chanx_right_in[97], chanx_right_in[139], chany_bottom_in[93], chanx_left_in[23], chanx_left_in[69], chanx_left_in[76], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size13_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_23_sram_inv[0:7]),
		.out(chany_top_out[93]));

	mux_2level_tapbuf_size13 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[34], chanx_right_in[87], chanx_right_in[101], chanx_right_in[140], chany_bottom_in[97], chanx_left_in[22], chanx_left_in[65], chanx_left_in[75], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size13_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_24_sram_inv[0:7]),
		.out(chany_top_out[97]));

	mux_2level_tapbuf_size13 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[35], chanx_right_in[88], chanx_right_in[105], chanx_right_in[142], chany_bottom_in[101], chanx_left_in[20], chanx_left_in[61], chanx_left_in[74], chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size13_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_25_sram_inv[0:7]),
		.out(chany_top_out[101]));

	mux_2level_tapbuf_size13 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[36], chanx_right_in[90], chanx_right_in[109], chanx_right_in[143], chany_bottom_in[105], chanx_left_in[19], chanx_left_in[57], chanx_left_in[72], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size13_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_26_sram_inv[0:7]),
		.out(chany_top_out[105]));

	mux_2level_tapbuf_size13 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[38], chanx_right_in[91], chanx_right_in[113], chanx_right_in[144], chany_bottom_in[109], chanx_left_in[18], chanx_left_in[53], chanx_left_in[71], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size13_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_27_sram_inv[0:7]),
		.out(chany_top_out[109]));

	mux_2level_tapbuf_size13 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[39], chanx_right_in[92], chanx_right_in[117], chanx_right_in[146], chany_bottom_in[113], chanx_left_in[16], chanx_left_in[49], chanx_left_in[70], chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size13_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_28_sram_inv[0:7]),
		.out(chany_top_out[113]));

	mux_2level_tapbuf_size13 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[40], chanx_right_in[94], chanx_right_in[121], chanx_right_in[147], chany_bottom_in[117], chanx_left_in[15], chanx_left_in[45], chanx_left_in[68], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size13_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_29_sram_inv[0:7]),
		.out(chany_top_out[117]));

	mux_2level_tapbuf_size13 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[42], chanx_right_in[95], chanx_right_in[125], chanx_right_in[148], chany_bottom_in[121], chanx_left_in[14], chanx_left_in[41], chanx_left_in[67], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size13_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_30_sram_inv[0:7]),
		.out(chany_top_out[121]));

	mux_2level_tapbuf_size13 mux_top_track_250 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[43], chanx_right_in[96], chanx_right_in[129], chanx_right_in[150], chany_bottom_in[125], chanx_left_in[12], chanx_left_in[37], chanx_left_in[66], chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size13_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_31_sram_inv[0:7]),
		.out(chany_top_out[125]));

	mux_2level_tapbuf_size13 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[44], chanx_right_in[98], chanx_right_in[133], chanx_right_in[151], chany_bottom_in[129], chanx_left_in[11], chanx_left_in[33], chanx_left_in[64], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size13_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_32_sram_inv[0:7]),
		.out(chany_top_out[129]));

	mux_2level_tapbuf_size13 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[46], chanx_right_in[99], chanx_right_in[137], chanx_right_in[152], chany_bottom_in[133], chanx_left_in[10], chanx_left_in[29], chanx_left_in[63], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size13_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_33_sram_inv[0:7]),
		.out(chany_top_out[133]));

	mux_2level_tapbuf_size13 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[47], chanx_right_in[100], chanx_right_in[141], chanx_right_in[154], chany_bottom_in[137], chanx_left_in[8], chanx_left_in[25], chanx_left_in[62], chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size13_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_34_sram_inv[0:7]),
		.out(chany_top_out[137]));

	mux_2level_tapbuf_size13 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[48], chanx_right_in[102], chanx_right_in[145], chanx_right_in[155], chany_bottom_in[141], chanx_left_in[7], chanx_left_in[21], chanx_left_in[60], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size13_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_35_sram_inv[0:7]),
		.out(chany_top_out[141]));

	mux_2level_tapbuf_size13 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[50], chanx_right_in[103], chanx_right_in[149], chanx_right_in[156], chany_bottom_in[145], chanx_left_in[6], chanx_left_in[17], chanx_left_in[59], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size13_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_36_sram_inv[0:7]),
		.out(chany_top_out[145]));

	mux_2level_tapbuf_size13 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[51], chanx_right_in[104], chanx_right_in[153], chanx_right_in[158], chany_bottom_in[149], chanx_left_in[4], chanx_left_in[13], chanx_left_in[58], chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size13_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_37_sram_inv[0:7]),
		.out(chany_top_out[149]));

	mux_2level_tapbuf_size13 mux_top_track_306 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[52], chanx_right_in[106], chanx_right_in[157], chanx_right_in[159], chany_bottom_in[153], chanx_left_in[3], chanx_left_in[9], chanx_left_in[56], chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size13_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_38_sram_inv[0:7]),
		.out(chany_top_out[153]));

	mux_2level_tapbuf_size13 mux_top_track_314 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[0:1], chanx_right_in[54], chanx_right_in[107], chany_bottom_in[157], chanx_left_in[2], chanx_left_in[5], chanx_left_in[55], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size13_39_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_39_sram_inv[0:7]),
		.out(chany_top_out[157]));

	mux_2level_tapbuf_size13 mux_left_track_3 (
		.in({chany_top_in[0:1], chany_top_in[54], chany_top_in[107], chanx_right_in[1], chany_bottom_in[52], chany_bottom_in[106], chany_bottom_in[157], chany_bottom_in[159], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_40_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_40_sram_inv[0:7]),
		.out(chanx_left_out[1]));

	mux_2level_tapbuf_size13 mux_left_track_11 (
		.in({chany_top_in[52], chany_top_in[106], chany_top_in[157], chany_top_in[159], chanx_right_in[5], chany_bottom_in[0:1], chany_bottom_in[54], chany_bottom_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_41_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_41_sram_inv[0:7]),
		.out(chanx_left_out[5]));

	mux_2level_tapbuf_size13 mux_left_track_19 (
		.in({chany_top_in[51], chany_top_in[104], chany_top_in[153], chany_top_in[158], chanx_right_in[9], chany_bottom_in[2], chany_bottom_in[5], chany_bottom_in[55], chany_bottom_in[108], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_42_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_42_sram_inv[0:7]),
		.out(chanx_left_out[9]));

	mux_2level_tapbuf_size13 mux_left_track_27 (
		.in({chany_top_in[50], chany_top_in[103], chany_top_in[149], chany_top_in[156], chanx_right_in[13], chany_bottom_in[3], chany_bottom_in[9], chany_bottom_in[56], chany_bottom_in[110], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_43_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_43_sram_inv[0:7]),
		.out(chanx_left_out[13]));

	mux_2level_tapbuf_size13 mux_left_track_35 (
		.in({chany_top_in[48], chany_top_in[102], chany_top_in[145], chany_top_in[155], chanx_right_in[17], chany_bottom_in[4], chany_bottom_in[13], chany_bottom_in[58], chany_bottom_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_44_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_44_sram_inv[0:7]),
		.out(chanx_left_out[17]));

	mux_2level_tapbuf_size13 mux_left_track_43 (
		.in({chany_top_in[47], chany_top_in[100], chany_top_in[141], chany_top_in[154], chanx_right_in[21], chany_bottom_in[6], chany_bottom_in[17], chany_bottom_in[59], chany_bottom_in[112], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_45_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_45_sram_inv[0:7]),
		.out(chanx_left_out[21]));

	mux_2level_tapbuf_size13 mux_left_track_51 (
		.in({chany_top_in[46], chany_top_in[99], chany_top_in[137], chany_top_in[152], chanx_right_in[25], chany_bottom_in[7], chany_bottom_in[21], chany_bottom_in[60], chany_bottom_in[114], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_46_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_46_sram_inv[0:7]),
		.out(chanx_left_out[25]));

	mux_2level_tapbuf_size13 mux_left_track_59 (
		.in({chany_top_in[44], chany_top_in[98], chany_top_in[133], chany_top_in[151], chanx_right_in[29], chany_bottom_in[8], chany_bottom_in[25], chany_bottom_in[62], chany_bottom_in[115], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size13_47_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_47_sram_inv[0:7]),
		.out(chanx_left_out[29]));

	mux_2level_tapbuf_size13 mux_left_track_67 (
		.in({chany_top_in[43], chany_top_in[96], chany_top_in[129], chany_top_in[150], chanx_right_in[33], chany_bottom_in[10], chany_bottom_in[29], chany_bottom_in[63], chany_bottom_in[116], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_48_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_48_sram_inv[0:7]),
		.out(chanx_left_out[33]));

	mux_2level_tapbuf_size13 mux_left_track_75 (
		.in({chany_top_in[42], chany_top_in[95], chany_top_in[125], chany_top_in[148], chanx_right_in[37], chany_bottom_in[11], chany_bottom_in[33], chany_bottom_in[64], chany_bottom_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_49_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_49_sram_inv[0:7]),
		.out(chanx_left_out[37]));

	mux_2level_tapbuf_size13 mux_left_track_83 (
		.in({chany_top_in[40], chany_top_in[94], chany_top_in[121], chany_top_in[147], chanx_right_in[41], chany_bottom_in[12], chany_bottom_in[37], chany_bottom_in[66], chany_bottom_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_50_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_50_sram_inv[0:7]),
		.out(chanx_left_out[41]));

	mux_2level_tapbuf_size13 mux_left_track_91 (
		.in({chany_top_in[39], chany_top_in[92], chany_top_in[117], chany_top_in[146], chanx_right_in[45], chany_bottom_in[14], chany_bottom_in[41], chany_bottom_in[67], chany_bottom_in[120], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_51_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_51_sram_inv[0:7]),
		.out(chanx_left_out[45]));

	mux_2level_tapbuf_size13 mux_left_track_99 (
		.in({chany_top_in[38], chany_top_in[91], chany_top_in[113], chany_top_in[144], chanx_right_in[49], chany_bottom_in[15], chany_bottom_in[45], chany_bottom_in[68], chany_bottom_in[122], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_52_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_52_sram_inv[0:7]),
		.out(chanx_left_out[49]));

	mux_2level_tapbuf_size13 mux_left_track_107 (
		.in({chany_top_in[36], chany_top_in[90], chany_top_in[109], chany_top_in[143], chanx_right_in[53], chany_bottom_in[16], chany_bottom_in[49], chany_bottom_in[70], chany_bottom_in[123], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_53_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_53_sram_inv[0:7]),
		.out(chanx_left_out[53]));

	mux_2level_tapbuf_size13 mux_left_track_115 (
		.in({chany_top_in[35], chany_top_in[88], chany_top_in[105], chany_top_in[142], chanx_right_in[57], chany_bottom_in[18], chany_bottom_in[53], chany_bottom_in[71], chany_bottom_in[124], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_54_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_54_sram_inv[0:7]),
		.out(chanx_left_out[57]));

	mux_2level_tapbuf_size13 mux_left_track_123 (
		.in({chany_top_in[34], chany_top_in[87], chany_top_in[101], chany_top_in[140], chanx_right_in[61], chany_bottom_in[19], chany_bottom_in[57], chany_bottom_in[72], chany_bottom_in[126], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_55_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_55_sram_inv[0:7]),
		.out(chanx_left_out[61]));

	mux_2level_tapbuf_size13 mux_left_track_131 (
		.in({chany_top_in[32], chany_top_in[86], chany_top_in[97], chany_top_in[139], chanx_right_in[65], chany_bottom_in[20], chany_bottom_in[61], chany_bottom_in[74], chany_bottom_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_56_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_56_sram_inv[0:7]),
		.out(chanx_left_out[65]));

	mux_2level_tapbuf_size13 mux_left_track_139 (
		.in({chany_top_in[31], chany_top_in[84], chany_top_in[93], chany_top_in[138], chanx_right_in[69], chany_bottom_in[22], chany_bottom_in[65], chany_bottom_in[75], chany_bottom_in[128], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_57_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_57_sram_inv[0:7]),
		.out(chanx_left_out[69]));

	mux_2level_tapbuf_size13 mux_left_track_147 (
		.in({chany_top_in[30], chany_top_in[83], chany_top_in[89], chany_top_in[136], chanx_right_in[73], chany_bottom_in[23], chany_bottom_in[69], chany_bottom_in[76], chany_bottom_in[130], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_58_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_58_sram_inv[0:7]),
		.out(chanx_left_out[73]));

	mux_2level_tapbuf_size13 mux_left_track_155 (
		.in({chany_top_in[28], chany_top_in[82], chany_top_in[85], chany_top_in[135], chanx_right_in[77], chany_bottom_in[24], chany_bottom_in[73], chany_bottom_in[78], chany_bottom_in[131], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_59_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_59_sram_inv[0:7]),
		.out(chanx_left_out[77]));

	mux_2level_tapbuf_size13 mux_left_track_163 (
		.in({chany_top_in[27], chany_top_in[80:81], chany_top_in[134], chanx_right_in[81], chany_bottom_in[26], chany_bottom_in[77], chany_bottom_in[79], chany_bottom_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_60_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_60_sram_inv[0:7]),
		.out(chanx_left_out[81]));

	mux_2level_tapbuf_size13 mux_left_track_171 (
		.in({chany_top_in[26], chany_top_in[77], chany_top_in[79], chany_top_in[132], chanx_right_in[85], chany_bottom_in[27], chany_bottom_in[80:81], chany_bottom_in[134], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_61_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_61_sram_inv[0:7]),
		.out(chanx_left_out[85]));

	mux_2level_tapbuf_size13 mux_left_track_179 (
		.in({chany_top_in[24], chany_top_in[73], chany_top_in[78], chany_top_in[131], chanx_right_in[89], chany_bottom_in[28], chany_bottom_in[82], chany_bottom_in[85], chany_bottom_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_62_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_62_sram_inv[0:7]),
		.out(chanx_left_out[89]));

	mux_2level_tapbuf_size13 mux_left_track_187 (
		.in({chany_top_in[23], chany_top_in[69], chany_top_in[76], chany_top_in[130], chanx_right_in[93], chany_bottom_in[30], chany_bottom_in[83], chany_bottom_in[89], chany_bottom_in[136], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size13_63_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_63_sram_inv[0:7]),
		.out(chanx_left_out[93]));

	mux_2level_tapbuf_size13 mux_left_track_195 (
		.in({chany_top_in[22], chany_top_in[65], chany_top_in[75], chany_top_in[128], chanx_right_in[97], chany_bottom_in[31], chany_bottom_in[84], chany_bottom_in[93], chany_bottom_in[138], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_64_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_64_sram_inv[0:7]),
		.out(chanx_left_out[97]));

	mux_2level_tapbuf_size13 mux_left_track_203 (
		.in({chany_top_in[20], chany_top_in[61], chany_top_in[74], chany_top_in[127], chanx_right_in[101], chany_bottom_in[32], chany_bottom_in[86], chany_bottom_in[97], chany_bottom_in[139], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_65_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_65_sram_inv[0:7]),
		.out(chanx_left_out[101]));

	mux_2level_tapbuf_size13 mux_left_track_211 (
		.in({chany_top_in[19], chany_top_in[57], chany_top_in[72], chany_top_in[126], chanx_right_in[105], chany_bottom_in[34], chany_bottom_in[87], chany_bottom_in[101], chany_bottom_in[140], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_66_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_66_sram_inv[0:7]),
		.out(chanx_left_out[105]));

	mux_2level_tapbuf_size13 mux_left_track_219 (
		.in({chany_top_in[18], chany_top_in[53], chany_top_in[71], chany_top_in[124], chanx_right_in[109], chany_bottom_in[35], chany_bottom_in[88], chany_bottom_in[105], chany_bottom_in[142], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_67_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_67_sram_inv[0:7]),
		.out(chanx_left_out[109]));

	mux_2level_tapbuf_size13 mux_left_track_227 (
		.in({chany_top_in[16], chany_top_in[49], chany_top_in[70], chany_top_in[123], chanx_right_in[113], chany_bottom_in[36], chany_bottom_in[90], chany_bottom_in[109], chany_bottom_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_68_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_68_sram_inv[0:7]),
		.out(chanx_left_out[113]));

	mux_2level_tapbuf_size13 mux_left_track_235 (
		.in({chany_top_in[15], chany_top_in[45], chany_top_in[68], chany_top_in[122], chanx_right_in[117], chany_bottom_in[38], chany_bottom_in[91], chany_bottom_in[113], chany_bottom_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_69_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_69_sram_inv[0:7]),
		.out(chanx_left_out[117]));

	mux_2level_tapbuf_size13 mux_left_track_243 (
		.in({chany_top_in[14], chany_top_in[41], chany_top_in[67], chany_top_in[120], chanx_right_in[121], chany_bottom_in[39], chany_bottom_in[92], chany_bottom_in[117], chany_bottom_in[146], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_70_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_70_sram_inv[0:7]),
		.out(chanx_left_out[121]));

	mux_2level_tapbuf_size13 mux_left_track_251 (
		.in({chany_top_in[12], chany_top_in[37], chany_top_in[66], chany_top_in[119], chanx_right_in[125], chany_bottom_in[40], chany_bottom_in[94], chany_bottom_in[121], chany_bottom_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_71_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_71_sram_inv[0:7]),
		.out(chanx_left_out[125]));

	mux_2level_tapbuf_size13 mux_left_track_259 (
		.in({chany_top_in[11], chany_top_in[33], chany_top_in[64], chany_top_in[118], chanx_right_in[129], chany_bottom_in[42], chany_bottom_in[95], chany_bottom_in[125], chany_bottom_in[148], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_72_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_72_sram_inv[0:7]),
		.out(chanx_left_out[129]));

	mux_2level_tapbuf_size13 mux_left_track_267 (
		.in({chany_top_in[10], chany_top_in[29], chany_top_in[63], chany_top_in[116], chanx_right_in[133], chany_bottom_in[43], chany_bottom_in[96], chany_bottom_in[129], chany_bottom_in[150], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_73_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_73_sram_inv[0:7]),
		.out(chanx_left_out[133]));

	mux_2level_tapbuf_size13 mux_left_track_275 (
		.in({chany_top_in[8], chany_top_in[25], chany_top_in[62], chany_top_in[115], chanx_right_in[137], chany_bottom_in[44], chany_bottom_in[98], chany_bottom_in[133], chany_bottom_in[151], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_74_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_74_sram_inv[0:7]),
		.out(chanx_left_out[137]));

	mux_2level_tapbuf_size13 mux_left_track_283 (
		.in({chany_top_in[7], chany_top_in[21], chany_top_in[60], chany_top_in[114], chanx_right_in[141], chany_bottom_in[46], chany_bottom_in[99], chany_bottom_in[137], chany_bottom_in[152], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_75_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_75_sram_inv[0:7]),
		.out(chanx_left_out[141]));

	mux_2level_tapbuf_size13 mux_left_track_291 (
		.in({chany_top_in[6], chany_top_in[17], chany_top_in[59], chany_top_in[112], chanx_right_in[145], chany_bottom_in[47], chany_bottom_in[100], chany_bottom_in[141], chany_bottom_in[154], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_76_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_76_sram_inv[0:7]),
		.out(chanx_left_out[145]));

	mux_2level_tapbuf_size13 mux_left_track_299 (
		.in({chany_top_in[4], chany_top_in[13], chany_top_in[58], chany_top_in[111], chanx_right_in[149], chany_bottom_in[48], chany_bottom_in[102], chany_bottom_in[145], chany_bottom_in[155], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_77_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_77_sram_inv[0:7]),
		.out(chanx_left_out[149]));

	mux_2level_tapbuf_size13 mux_left_track_307 (
		.in({chany_top_in[3], chany_top_in[9], chany_top_in[56], chany_top_in[110], chanx_right_in[153], chany_bottom_in[50], chany_bottom_in[103], chany_bottom_in[149], chany_bottom_in[156], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_78_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_78_sram_inv[0:7]),
		.out(chanx_left_out[153]));

	mux_2level_tapbuf_size13 mux_left_track_315 (
		.in({chany_top_in[2], chany_top_in[5], chany_top_in[55], chany_top_in[108], chanx_right_in[157], chany_bottom_in[51], chany_bottom_in[104], chany_bottom_in[153], chany_bottom_in[158], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size13_79_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_79_sram_inv[0:7]),
		.out(chanx_left_out[157]));

	mux_2level_tapbuf_size13_mem mem_top_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_0_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_1_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_2_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_3_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_4_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_5_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_6_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_7_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_8_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_9_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_10_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_11_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_12_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_13_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_14_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_15_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_16_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_17_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_18_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_19_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_20_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_21_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_22_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_23_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_24_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_25_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_26_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_27_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_28_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_29_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_30_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_31_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_32_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_33_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_34_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_35_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_36_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_37_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_38_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_39_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_39_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_3 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size42_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_40_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_40_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_11 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_41_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_41_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_19 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_42_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_42_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_27 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_43_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_43_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_35 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_44_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_44_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_43 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_45_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_45_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_51 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_46_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_46_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_59 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_47_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_47_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_67 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_48_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_48_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_75 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_49_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_49_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_83 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_50_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_50_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_91 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_51_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_51_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_99 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_52_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_52_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_107 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_53_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_53_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_115 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_54_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_54_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_123 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_55_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_55_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_131 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_56_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_56_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_139 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_57_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_57_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_147 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_58_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_58_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_155 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_59_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_59_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_163 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_60_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_60_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_171 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_61_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_61_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_179 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_62_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_62_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_187 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_63_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_63_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_195 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_64_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_64_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_203 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_65_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_65_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_211 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_66_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_66_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_219 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_67_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_67_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_227 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_68_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_68_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_235 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_69_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_69_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_243 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_70_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_70_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_251 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_71_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_71_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_259 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_72_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_72_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_267 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_73_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_73_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_275 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_74_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_74_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_283 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_75_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_75_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_291 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_76_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_76_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_299 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_77_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_77_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_307 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_78_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_78_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_315 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_78_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_79_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_79_sram_inv[0:7]));

	mux_2level_tapbuf_size29 mux_right_track_2 (
		.in({chany_top_in[52], chany_top_in[106], chany_top_in[157], chany_top_in[159], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[51], chany_bottom_in[104], chany_bottom_in[153], chany_bottom_in[158], chanx_left_in[1]}),
		.sram(mux_2level_tapbuf_size29_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_0_sram_inv[0:11]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size29_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_0_sram_inv[0:11]));

	mux_2level_tapbuf_size27 mux_right_track_10 (
		.in({chany_top_in[0:1], chany_top_in[54], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[50], chany_bottom_in[149], chanx_left_in[5]}),
		.sram(mux_2level_tapbuf_size27_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_0_sram_inv[0:11]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size27 mux_right_track_18 (
		.in({chany_top_in[2], chany_top_in[5], chany_top_in[55], chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[48], chany_bottom_in[145], chanx_left_in[9]}),
		.sram(mux_2level_tapbuf_size27_1_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_1_sram_inv[0:11]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size27 mux_right_track_26 (
		.in({chany_top_in[3], chany_top_in[9], chany_top_in[56], chany_top_in[110], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[47], chany_bottom_in[141], chanx_left_in[13]}),
		.sram(mux_2level_tapbuf_size27_2_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_2_sram_inv[0:11]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size27 mux_right_track_34 (
		.in({chany_top_in[4], chany_top_in[13], chany_top_in[58], chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[46], chany_bottom_in[137], chanx_left_in[17]}),
		.sram(mux_2level_tapbuf_size27_3_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_3_sram_inv[0:11]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size27 mux_right_track_42 (
		.in({chany_top_in[6], chany_top_in[17], chany_top_in[59], chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[44], chany_bottom_in[133], chanx_left_in[21]}),
		.sram(mux_2level_tapbuf_size27_4_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_4_sram_inv[0:11]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size27 mux_right_track_50 (
		.in({chany_top_in[7], chany_top_in[21], chany_top_in[60], chany_top_in[114], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[43], chany_bottom_in[129], chanx_left_in[25]}),
		.sram(mux_2level_tapbuf_size27_5_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_5_sram_inv[0:11]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size27 mux_right_track_58 (
		.in({chany_top_in[8], chany_top_in[25], chany_top_in[62], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[42], chany_bottom_in[125], chanx_left_in[29]}),
		.sram(mux_2level_tapbuf_size27_6_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size27_6_sram_inv[0:11]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size27_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_0_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_1_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_1_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_2_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_2_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_3_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_3_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_4_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_4_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_5_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_5_sram_inv[0:11]));

	mux_2level_tapbuf_size27_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size27_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size27_6_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size27_6_sram_inv[0:11]));

	mux_2level_tapbuf_size26 mux_right_track_66 (
		.in({chany_top_in[10], chany_top_in[29], chany_top_in[63], chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[40], chany_bottom_in[121], chanx_left_in[33]}),
		.sram(mux_2level_tapbuf_size26_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_0_sram_inv[0:11]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size26 mux_right_track_74 (
		.in({chany_top_in[11], chany_top_in[33], chany_top_in[64], chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[39], chany_bottom_in[117], chanx_left_in[37]}),
		.sram(mux_2level_tapbuf_size26_1_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_1_sram_inv[0:11]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size26 mux_right_track_82 (
		.in({chany_top_in[12], chany_top_in[37], chany_top_in[66], chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[38], chany_bottom_in[113], chanx_left_in[41]}),
		.sram(mux_2level_tapbuf_size26_2_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_2_sram_inv[0:11]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size26 mux_right_track_90 (
		.in({chany_top_in[14], chany_top_in[41], chany_top_in[67], chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[36], chany_bottom_in[109], chanx_left_in[45]}),
		.sram(mux_2level_tapbuf_size26_3_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_3_sram_inv[0:11]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size26 mux_right_track_98 (
		.in({chany_top_in[15], chany_top_in[45], chany_top_in[68], chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[35], chany_bottom_in[105], chanx_left_in[49]}),
		.sram(mux_2level_tapbuf_size26_4_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_4_sram_inv[0:11]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size26 mux_right_track_106 (
		.in({chany_top_in[16], chany_top_in[49], chany_top_in[70], chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[34], chany_bottom_in[101], chanx_left_in[53]}),
		.sram(mux_2level_tapbuf_size26_5_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_5_sram_inv[0:11]),
		.out(chanx_right_out[53]));

	mux_2level_tapbuf_size26 mux_right_track_114 (
		.in({chany_top_in[18], chany_top_in[53], chany_top_in[71], chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[32], chany_bottom_in[97], chanx_left_in[57]}),
		.sram(mux_2level_tapbuf_size26_6_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_6_sram_inv[0:11]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size26 mux_right_track_122 (
		.in({chany_top_in[19], chany_top_in[57], chany_top_in[72], chany_top_in[126], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[31], chany_bottom_in[93], chanx_left_in[61]}),
		.sram(mux_2level_tapbuf_size26_7_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_7_sram_inv[0:11]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size26 mux_right_track_130 (
		.in({chany_top_in[20], chany_top_in[61], chany_top_in[74], chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[30], chany_bottom_in[89], chanx_left_in[65]}),
		.sram(mux_2level_tapbuf_size26_8_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_8_sram_inv[0:11]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size26 mux_right_track_138 (
		.in({chany_top_in[22], chany_top_in[65], chany_top_in[75], chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[28], chany_bottom_in[85], chanx_left_in[69]}),
		.sram(mux_2level_tapbuf_size26_9_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_9_sram_inv[0:11]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size26 mux_right_track_146 (
		.in({chany_top_in[23], chany_top_in[69], chany_top_in[76], chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[27], chany_bottom_in[81], chanx_left_in[73]}),
		.sram(mux_2level_tapbuf_size26_10_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_10_sram_inv[0:11]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size26 mux_right_track_154 (
		.in({chany_top_in[24], chany_top_in[73], chany_top_in[78], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[26], chany_bottom_in[77], chanx_left_in[77]}),
		.sram(mux_2level_tapbuf_size26_11_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_11_sram_inv[0:11]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size26 mux_right_track_162 (
		.in({chany_top_in[26], chany_top_in[77], chany_top_in[79], chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[24], chany_bottom_in[73], chanx_left_in[81]}),
		.sram(mux_2level_tapbuf_size26_12_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_12_sram_inv[0:11]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size26 mux_right_track_170 (
		.in({chany_top_in[27], chany_top_in[80:81], chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[23], chany_bottom_in[69], chanx_left_in[85]}),
		.sram(mux_2level_tapbuf_size26_13_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_13_sram_inv[0:11]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size26 mux_right_track_178 (
		.in({chany_top_in[28], chany_top_in[82], chany_top_in[85], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[22], chany_bottom_in[65], chanx_left_in[89]}),
		.sram(mux_2level_tapbuf_size26_14_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_14_sram_inv[0:11]),
		.out(chanx_right_out[89]));

	mux_2level_tapbuf_size26 mux_right_track_186 (
		.in({chany_top_in[30], chany_top_in[83], chany_top_in[89], chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[20], chany_bottom_in[61], chanx_left_in[93]}),
		.sram(mux_2level_tapbuf_size26_15_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_15_sram_inv[0:11]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size26 mux_right_track_194 (
		.in({chany_top_in[31], chany_top_in[84], chany_top_in[93], chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[19], chany_bottom_in[57], chanx_left_in[97]}),
		.sram(mux_2level_tapbuf_size26_16_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_16_sram_inv[0:11]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size26 mux_right_track_202 (
		.in({chany_top_in[32], chany_top_in[86], chany_top_in[97], chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[18], chany_bottom_in[53], chanx_left_in[101]}),
		.sram(mux_2level_tapbuf_size26_17_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_17_sram_inv[0:11]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size26 mux_right_track_210 (
		.in({chany_top_in[34], chany_top_in[87], chany_top_in[101], chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[16], chany_bottom_in[49], chanx_left_in[105]}),
		.sram(mux_2level_tapbuf_size26_18_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_18_sram_inv[0:11]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size26 mux_right_track_218 (
		.in({chany_top_in[35], chany_top_in[88], chany_top_in[105], chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[15], chany_bottom_in[45], chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size26_19_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_19_sram_inv[0:11]),
		.out(chanx_right_out[109]));

	mux_2level_tapbuf_size26 mux_right_track_226 (
		.in({chany_top_in[36], chany_top_in[90], chany_top_in[109], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[14], chany_bottom_in[41], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size26_20_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_20_sram_inv[0:11]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size26 mux_right_track_234 (
		.in({chany_top_in[38], chany_top_in[91], chany_top_in[113], chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[12], chany_bottom_in[37], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size26_21_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_21_sram_inv[0:11]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size26 mux_right_track_242 (
		.in({chany_top_in[39], chany_top_in[92], chany_top_in[117], chany_top_in[146], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[11], chany_bottom_in[33], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size26_22_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_22_sram_inv[0:11]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size26 mux_right_track_250 (
		.in({chany_top_in[40], chany_top_in[94], chany_top_in[121], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[10], chany_bottom_in[29], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size26_23_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_23_sram_inv[0:11]),
		.out(chanx_right_out[125]));

	mux_2level_tapbuf_size26 mux_right_track_258 (
		.in({chany_top_in[42], chany_top_in[95], chany_top_in[125], chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[8], chany_bottom_in[25], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size26_24_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_24_sram_inv[0:11]),
		.out(chanx_right_out[129]));

	mux_2level_tapbuf_size26 mux_right_track_266 (
		.in({chany_top_in[43], chany_top_in[96], chany_top_in[129], chany_top_in[150], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[7], chany_bottom_in[21], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size26_25_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_25_sram_inv[0:11]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size26 mux_right_track_274 (
		.in({chany_top_in[44], chany_top_in[98], chany_top_in[133], chany_top_in[151], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[6], chany_bottom_in[17], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size26_26_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_26_sram_inv[0:11]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size26 mux_right_track_282 (
		.in({chany_top_in[46], chany_top_in[99], chany_top_in[137], chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[4], chany_bottom_in[13], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size26_27_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_27_sram_inv[0:11]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size26 mux_right_track_290 (
		.in({chany_top_in[47], chany_top_in[100], chany_top_in[141], chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[3], chany_bottom_in[9], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size26_28_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_28_sram_inv[0:11]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size26 mux_right_track_298 (
		.in({chany_top_in[48], chany_top_in[102], chany_top_in[145], chany_top_in[155], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[2], chany_bottom_in[5], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size26_29_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_29_sram_inv[0:11]),
		.out(chanx_right_out[149]));

	mux_2level_tapbuf_size26 mux_right_track_306 (
		.in({chany_top_in[50], chany_top_in[103], chany_top_in[149], chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[0:1], chanx_left_in[153]}),
		.sram(mux_2level_tapbuf_size26_30_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size26_30_sram_inv[0:11]),
		.out(chanx_right_out[153]));

	mux_2level_tapbuf_size26_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size27_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_0_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_1_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_1_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_2_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_2_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_3_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_3_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_4_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_4_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_5_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_5_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_6_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_6_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_7_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_7_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_8_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_8_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_9_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_9_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_10_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_10_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_11_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_11_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_12_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_12_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_13_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_13_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_14_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_14_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_15_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_15_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_16_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_16_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_17_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_17_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_18_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_18_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_19_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_19_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_20_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_20_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_21_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_21_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_22_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_22_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_23_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_23_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_24_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_24_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_25_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_25_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_26_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_26_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_27_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_27_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_28_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_28_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_29_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_29_sram_inv[0:11]));

	mux_2level_tapbuf_size26_mem mem_right_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size26_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size26_30_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size26_30_sram_inv[0:11]));

	mux_2level_tapbuf_size25 mux_right_track_314 (
		.in({chany_top_in[51], chany_top_in[104], chany_top_in[153], chany_top_in[158], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[157], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size25_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size25_0_sram_inv[0:11]),
		.out(chanx_right_out[157]));

	mux_2level_tapbuf_size25_mem mem_right_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size26_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size25_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size25_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size25_0_sram_inv[0:11]));

	mux_2level_tapbuf_size46 mux_bottom_track_3 (
		.in({chany_top_in[1], chanx_right_in[51], chanx_right_in[104], chanx_right_in[153], chanx_right_in[158], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[2], chanx_left_in[5], chanx_left_in[55], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size46_0_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size46_0_sram_inv[0:13]),
		.out(chany_bottom_out[1]));

	mux_2level_tapbuf_size46_mem mem_bottom_track_3 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size25_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size46_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size46_0_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size46_0_sram_inv[0:13]));

	mux_2level_tapbuf_size44 mux_bottom_track_11 (
		.in({chany_top_in[5], chanx_right_in[50], chanx_right_in[149], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[3], chanx_left_in[9], chanx_left_in[56], chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size44_0_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_0_sram_inv[0:13]),
		.out(chany_bottom_out[5]));

	mux_2level_tapbuf_size44 mux_bottom_track_19 (
		.in({chany_top_in[9], chanx_right_in[48], chanx_right_in[145], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[4], chanx_left_in[13], chanx_left_in[58], chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size44_1_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_1_sram_inv[0:13]),
		.out(chany_bottom_out[9]));

	mux_2level_tapbuf_size44 mux_bottom_track_27 (
		.in({chany_top_in[13], chanx_right_in[47], chanx_right_in[141], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[6], chanx_left_in[17], chanx_left_in[59], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size44_2_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_2_sram_inv[0:13]),
		.out(chany_bottom_out[13]));

	mux_2level_tapbuf_size44 mux_bottom_track_35 (
		.in({chany_top_in[17], chanx_right_in[46], chanx_right_in[137], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[7], chanx_left_in[21], chanx_left_in[60], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size44_3_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_3_sram_inv[0:13]),
		.out(chany_bottom_out[17]));

	mux_2level_tapbuf_size44 mux_bottom_track_43 (
		.in({chany_top_in[21], chanx_right_in[44], chanx_right_in[133], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[8], chanx_left_in[25], chanx_left_in[62], chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size44_4_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_4_sram_inv[0:13]),
		.out(chany_bottom_out[21]));

	mux_2level_tapbuf_size44 mux_bottom_track_51 (
		.in({chany_top_in[25], chanx_right_in[43], chanx_right_in[129], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[10], chanx_left_in[29], chanx_left_in[63], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size44_5_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_5_sram_inv[0:13]),
		.out(chany_bottom_out[25]));

	mux_2level_tapbuf_size44 mux_bottom_track_59 (
		.in({chany_top_in[29], chanx_right_in[42], chanx_right_in[125], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[11], chanx_left_in[33], chanx_left_in[64], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size44_6_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_6_sram_inv[0:13]),
		.out(chany_bottom_out[29]));

	mux_2level_tapbuf_size44 mux_bottom_track_67 (
		.in({chany_top_in[33], chanx_right_in[40], chanx_right_in[121], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[12], chanx_left_in[37], chanx_left_in[66], chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size44_7_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_7_sram_inv[0:13]),
		.out(chany_bottom_out[33]));

	mux_2level_tapbuf_size44 mux_bottom_track_75 (
		.in({chany_top_in[37], chanx_right_in[39], chanx_right_in[117], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[14], chanx_left_in[41], chanx_left_in[67], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size44_8_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_8_sram_inv[0:13]),
		.out(chany_bottom_out[37]));

	mux_2level_tapbuf_size44 mux_bottom_track_83 (
		.in({chany_top_in[41], chanx_right_in[38], chanx_right_in[113], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[15], chanx_left_in[45], chanx_left_in[68], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size44_9_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_9_sram_inv[0:13]),
		.out(chany_bottom_out[41]));

	mux_2level_tapbuf_size44 mux_bottom_track_91 (
		.in({chany_top_in[45], chanx_right_in[36], chanx_right_in[109], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[16], chanx_left_in[49], chanx_left_in[70], chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size44_10_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_10_sram_inv[0:13]),
		.out(chany_bottom_out[45]));

	mux_2level_tapbuf_size44 mux_bottom_track_99 (
		.in({chany_top_in[49], chanx_right_in[35], chanx_right_in[105], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[18], chanx_left_in[53], chanx_left_in[71], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size44_11_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_11_sram_inv[0:13]),
		.out(chany_bottom_out[49]));

	mux_2level_tapbuf_size44 mux_bottom_track_107 (
		.in({chany_top_in[53], chanx_right_in[34], chanx_right_in[101], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[19], chanx_left_in[57], chanx_left_in[72], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size44_12_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_12_sram_inv[0:13]),
		.out(chany_bottom_out[53]));

	mux_2level_tapbuf_size44 mux_bottom_track_115 (
		.in({chany_top_in[57], chanx_right_in[32], chanx_right_in[97], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[20], chanx_left_in[61], chanx_left_in[74], chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size44_13_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_13_sram_inv[0:13]),
		.out(chany_bottom_out[57]));

	mux_2level_tapbuf_size44 mux_bottom_track_123 (
		.in({chany_top_in[61], chanx_right_in[31], chanx_right_in[93], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[22], chanx_left_in[65], chanx_left_in[75], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size44_14_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size44_14_sram_inv[0:13]),
		.out(chany_bottom_out[61]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_11 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size46_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_0_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_0_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_19 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_1_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_1_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_27 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_2_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_2_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_35 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_3_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_3_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_43 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_4_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_4_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_51 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_5_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_5_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_59 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_6_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_6_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_67 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_7_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_7_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_75 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_8_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_8_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_83 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_9_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_9_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_91 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_10_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_10_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_99 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_11_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_11_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_107 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_12_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_12_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_115 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_13_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_13_sram_inv[0:13]));

	mux_2level_tapbuf_size44_mem mem_bottom_track_123 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size44_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size44_14_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size44_14_sram_inv[0:13]));

	mux_2level_tapbuf_size43 mux_bottom_track_131 (
		.in({chany_top_in[65], chanx_right_in[30], chanx_right_in[89], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[23], chanx_left_in[69], chanx_left_in[76], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size43_0_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_0_sram_inv[0:13]),
		.out(chany_bottom_out[65]));

	mux_2level_tapbuf_size43 mux_bottom_track_139 (
		.in({chany_top_in[69], chanx_right_in[28], chanx_right_in[85], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[24], chanx_left_in[73], chanx_left_in[78], chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size43_1_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_1_sram_inv[0:13]),
		.out(chany_bottom_out[69]));

	mux_2level_tapbuf_size43 mux_bottom_track_147 (
		.in({chany_top_in[73], chanx_right_in[27], chanx_right_in[81], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[26], chanx_left_in[77], chanx_left_in[79], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size43_2_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_2_sram_inv[0:13]),
		.out(chany_bottom_out[73]));

	mux_2level_tapbuf_size43 mux_bottom_track_155 (
		.in({chany_top_in[77], chanx_right_in[26], chanx_right_in[77], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[27], chanx_left_in[80:81], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size43_3_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_3_sram_inv[0:13]),
		.out(chany_bottom_out[77]));

	mux_2level_tapbuf_size43 mux_bottom_track_163 (
		.in({chany_top_in[81], chanx_right_in[24], chanx_right_in[73], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[28], chanx_left_in[82], chanx_left_in[85], chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size43_4_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_4_sram_inv[0:13]),
		.out(chany_bottom_out[81]));

	mux_2level_tapbuf_size43 mux_bottom_track_171 (
		.in({chany_top_in[85], chanx_right_in[23], chanx_right_in[69], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[30], chanx_left_in[83], chanx_left_in[89], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size43_5_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_5_sram_inv[0:13]),
		.out(chany_bottom_out[85]));

	mux_2level_tapbuf_size43 mux_bottom_track_179 (
		.in({chany_top_in[89], chanx_right_in[22], chanx_right_in[65], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[31], chanx_left_in[84], chanx_left_in[93], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size43_6_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_6_sram_inv[0:13]),
		.out(chany_bottom_out[89]));

	mux_2level_tapbuf_size43 mux_bottom_track_187 (
		.in({chany_top_in[93], chanx_right_in[20], chanx_right_in[61], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[32], chanx_left_in[86], chanx_left_in[97], chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size43_7_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_7_sram_inv[0:13]),
		.out(chany_bottom_out[93]));

	mux_2level_tapbuf_size43 mux_bottom_track_195 (
		.in({chany_top_in[97], chanx_right_in[19], chanx_right_in[57], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[34], chanx_left_in[87], chanx_left_in[101], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size43_8_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_8_sram_inv[0:13]),
		.out(chany_bottom_out[97]));

	mux_2level_tapbuf_size43 mux_bottom_track_203 (
		.in({chany_top_in[101], chanx_right_in[18], chanx_right_in[53], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[35], chanx_left_in[88], chanx_left_in[105], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size43_9_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_9_sram_inv[0:13]),
		.out(chany_bottom_out[101]));

	mux_2level_tapbuf_size43 mux_bottom_track_211 (
		.in({chany_top_in[105], chanx_right_in[16], chanx_right_in[49], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[36], chanx_left_in[90], chanx_left_in[109], chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size43_10_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_10_sram_inv[0:13]),
		.out(chany_bottom_out[105]));

	mux_2level_tapbuf_size43 mux_bottom_track_219 (
		.in({chany_top_in[109], chanx_right_in[15], chanx_right_in[45], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[38], chanx_left_in[91], chanx_left_in[113], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size43_11_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_11_sram_inv[0:13]),
		.out(chany_bottom_out[109]));

	mux_2level_tapbuf_size43 mux_bottom_track_227 (
		.in({chany_top_in[113], chanx_right_in[14], chanx_right_in[41], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[39], chanx_left_in[92], chanx_left_in[117], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size43_12_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_12_sram_inv[0:13]),
		.out(chany_bottom_out[113]));

	mux_2level_tapbuf_size43 mux_bottom_track_235 (
		.in({chany_top_in[117], chanx_right_in[12], chanx_right_in[37], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[40], chanx_left_in[94], chanx_left_in[121], chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size43_13_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_13_sram_inv[0:13]),
		.out(chany_bottom_out[117]));

	mux_2level_tapbuf_size43 mux_bottom_track_243 (
		.in({chany_top_in[121], chanx_right_in[11], chanx_right_in[33], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[42], chanx_left_in[95], chanx_left_in[125], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size43_14_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_14_sram_inv[0:13]),
		.out(chany_bottom_out[121]));

	mux_2level_tapbuf_size43 mux_bottom_track_251 (
		.in({chany_top_in[125], chanx_right_in[10], chanx_right_in[29], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[43], chanx_left_in[96], chanx_left_in[129], chanx_left_in[150]}),
		.sram(mux_2level_tapbuf_size43_15_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_15_sram_inv[0:13]),
		.out(chany_bottom_out[125]));

	mux_2level_tapbuf_size43 mux_bottom_track_259 (
		.in({chany_top_in[129], chanx_right_in[8], chanx_right_in[25], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[44], chanx_left_in[98], chanx_left_in[133], chanx_left_in[151]}),
		.sram(mux_2level_tapbuf_size43_16_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_16_sram_inv[0:13]),
		.out(chany_bottom_out[129]));

	mux_2level_tapbuf_size43 mux_bottom_track_267 (
		.in({chany_top_in[133], chanx_right_in[7], chanx_right_in[21], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[46], chanx_left_in[99], chanx_left_in[137], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size43_17_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_17_sram_inv[0:13]),
		.out(chany_bottom_out[133]));

	mux_2level_tapbuf_size43 mux_bottom_track_275 (
		.in({chany_top_in[137], chanx_right_in[6], chanx_right_in[17], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[47], chanx_left_in[100], chanx_left_in[141], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size43_18_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_18_sram_inv[0:13]),
		.out(chany_bottom_out[137]));

	mux_2level_tapbuf_size43 mux_bottom_track_283 (
		.in({chany_top_in[141], chanx_right_in[4], chanx_right_in[13], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[48], chanx_left_in[102], chanx_left_in[145], chanx_left_in[155]}),
		.sram(mux_2level_tapbuf_size43_19_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_19_sram_inv[0:13]),
		.out(chany_bottom_out[141]));

	mux_2level_tapbuf_size43 mux_bottom_track_291 (
		.in({chany_top_in[145], chanx_right_in[3], chanx_right_in[9], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[50], chanx_left_in[103], chanx_left_in[149], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size43_20_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_20_sram_inv[0:13]),
		.out(chany_bottom_out[145]));

	mux_2level_tapbuf_size43 mux_bottom_track_299 (
		.in({chany_top_in[149], chanx_right_in[2], chanx_right_in[5], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[51], chanx_left_in[104], chanx_left_in[153], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size43_21_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_21_sram_inv[0:13]),
		.out(chany_bottom_out[149]));

	mux_2level_tapbuf_size43 mux_bottom_track_307 (
		.in({chany_top_in[153], chanx_right_in[0:1], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[52], chanx_left_in[106], chanx_left_in[157], chanx_left_in[159]}),
		.sram(mux_2level_tapbuf_size43_22_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size43_22_sram_inv[0:13]),
		.out(chany_bottom_out[153]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_131 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size44_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_0_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_0_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_139 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_1_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_1_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_147 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_2_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_2_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_155 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_3_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_3_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_163 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_4_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_4_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_171 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_5_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_5_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_179 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_6_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_6_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_187 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_7_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_7_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_195 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_8_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_8_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_203 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_9_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_9_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_211 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_10_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_10_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_219 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_11_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_11_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_227 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_12_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_12_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_235 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_13_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_13_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_243 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_14_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_14_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_251 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_15_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_15_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_259 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_16_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_16_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_267 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_17_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_17_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_275 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_18_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_18_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_283 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_19_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_19_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_291 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_20_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_20_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_299 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_21_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_21_sram_inv[0:13]));

	mux_2level_tapbuf_size43_mem mem_bottom_track_307 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size43_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size43_22_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size43_22_sram_inv[0:13]));

	mux_2level_tapbuf_size42 mux_bottom_track_315 (
		.in({chany_top_in[157], chanx_right_in[157], bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[0:1], chanx_left_in[54], chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size42_0_sram[0:13]),
		.sram_inv(mux_2level_tapbuf_size42_0_sram_inv[0:13]),
		.out(chany_bottom_out[157]));

	mux_2level_tapbuf_size42_mem mem_bottom_track_315 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size43_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size42_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size42_0_sram[0:13]),
		.mem_outb(mux_2level_tapbuf_size42_0_sram_inv[0:13]));

endmodule
// ----- END Verilog module for sb_1__4_ -----

//----- Default net type -----
`default_nettype wire



