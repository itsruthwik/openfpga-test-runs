//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[4][3]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug 20 23:36:48 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_4__3_ -----
module sb_4__3_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_,
                chanx_right_in,
                chany_bottom_in,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:41] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_;
//----- INPUT PORTS -----
input [0:41] chanx_right_in;
//----- INPUT PORTS -----
input [0:41] chany_bottom_in;
//----- INPUT PORTS -----
input [0:41] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:41] chany_top_out;
//----- OUTPUT PORTS -----
output [0:41] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:41] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:41] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:9] mux_2level_tapbuf_size20_0_sram;
wire [0:9] mux_2level_tapbuf_size20_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size20_mem_0_ccff_tail;
wire [0:9] mux_2level_tapbuf_size21_0_sram;
wire [0:9] mux_2level_tapbuf_size21_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size21_1_sram;
wire [0:9] mux_2level_tapbuf_size21_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size21_mem_0_ccff_tail;
wire [0:9] mux_2level_tapbuf_size22_0_sram;
wire [0:9] mux_2level_tapbuf_size22_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_1_sram;
wire [0:9] mux_2level_tapbuf_size22_1_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_2_sram;
wire [0:9] mux_2level_tapbuf_size22_2_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_3_sram;
wire [0:9] mux_2level_tapbuf_size22_3_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_4_sram;
wire [0:9] mux_2level_tapbuf_size22_4_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_5_sram;
wire [0:9] mux_2level_tapbuf_size22_5_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_6_sram;
wire [0:9] mux_2level_tapbuf_size22_6_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_7_sram;
wire [0:9] mux_2level_tapbuf_size22_7_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_8_sram;
wire [0:9] mux_2level_tapbuf_size22_8_sram_inv;
wire [0:9] mux_2level_tapbuf_size22_9_sram;
wire [0:9] mux_2level_tapbuf_size22_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size22_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size22_mem_9_ccff_tail;
wire [0:9] mux_2level_tapbuf_size23_0_sram;
wire [0:9] mux_2level_tapbuf_size23_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_1_sram;
wire [0:9] mux_2level_tapbuf_size23_1_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_2_sram;
wire [0:9] mux_2level_tapbuf_size23_2_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_3_sram;
wire [0:9] mux_2level_tapbuf_size23_3_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_4_sram;
wire [0:9] mux_2level_tapbuf_size23_4_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_5_sram;
wire [0:9] mux_2level_tapbuf_size23_5_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_6_sram;
wire [0:9] mux_2level_tapbuf_size23_6_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_7_sram;
wire [0:9] mux_2level_tapbuf_size23_7_sram_inv;
wire [0:9] mux_2level_tapbuf_size23_8_sram;
wire [0:9] mux_2level_tapbuf_size23_8_sram_inv;
wire [0:0] mux_2level_tapbuf_size23_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size23_mem_8_ccff_tail;
wire [0:5] mux_2level_tapbuf_size6_0_sram;
wire [0:5] mux_2level_tapbuf_size6_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_1_sram;
wire [0:5] mux_2level_tapbuf_size6_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_1_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size23 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[16], chanx_right_in[30], chanx_left_in[0], chanx_left_in[3], chanx_left_in[14], chanx_left_in[29]}),
		.sram(mux_2level_tapbuf_size23_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_0_sram_inv[0:9]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size23 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[8], chanx_right_in[22], chanx_right_in[27], chanx_right_in[37], chanx_left_in[8], chanx_left_in[22], chanx_left_in[27], chanx_left_in[37]}),
		.sram(mux_2level_tapbuf_size23_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_1_sram_inv[0:9]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size23 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[9], chanx_right_in[24], chanx_right_in[31], chanx_right_in[38], chanx_left_in[6], chanx_left_in[21], chanx_left_in[23], chanx_left_in[36]}),
		.sram(mux_2level_tapbuf_size23_2_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_2_sram_inv[0:9]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size23 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[10], chanx_right_in[25], chanx_right_in[35], chanx_right_in[40], chanx_left_in[5], chanx_left_in[19:20], chanx_left_in[34]}),
		.sram(mux_2level_tapbuf_size23_3_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_3_sram_inv[0:9]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size23 mux_left_track_25 (
		.in({chany_top_in[10], chany_top_in[25], chany_top_in[35], chany_top_in[40], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[17], chany_bottom_in[32], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_}),
		.sram(mux_2level_tapbuf_size23_4_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_4_sram_inv[0:9]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size23 mux_left_track_41 (
		.in({chany_top_in[8], chany_top_in[22], chany_top_in[27], chany_top_in[37], chany_bottom_in[5], chany_bottom_in[19:20], chany_bottom_in[34], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size23_5_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_5_sram_inv[0:9]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size23 mux_left_track_49 (
		.in({chany_top_in[6], chany_top_in[21], chany_top_in[23], chany_top_in[36], chany_bottom_in[6], chany_bottom_in[21], chany_bottom_in[23], chany_bottom_in[36], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_}),
		.sram(mux_2level_tapbuf_size23_6_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_6_sram_inv[0:9]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size23 mux_left_track_57 (
		.in({chany_top_in[5], chany_top_in[19:20], chany_top_in[34], chany_bottom_in[8], chany_bottom_in[22], chany_bottom_in[27], chany_bottom_in[37], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_}),
		.sram(mux_2level_tapbuf_size23_7_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_7_sram_inv[0:9]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size23 mux_left_track_65 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[18], chany_top_in[33], chany_bottom_in[9], chany_bottom_in[24], chany_bottom_in[31], chany_bottom_in[38], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_}),
		.sram(mux_2level_tapbuf_size23_8_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size23_8_sram_inv[0:9]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size23_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size23_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_0_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_1_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_2_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_2_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_3_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_3_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_4_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_4_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_5_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_5_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_6_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_6_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_7_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_7_sram_inv[0:9]));

	mux_2level_tapbuf_size23_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size23_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size23_8_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size23_8_sram_inv[0:9]));

	mux_2level_tapbuf_size22 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[17], chanx_right_in[32], chanx_left_in[13], chanx_left_in[28], chanx_left_in[41]}),
		.sram(mux_2level_tapbuf_size22_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_0_sram_inv[0:9]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size22 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[4], chanx_right_in[15], chanx_right_in[18], chanx_right_in[33], chanx_left_in[12], chanx_left_in[26], chanx_left_in[39]}),
		.sram(mux_2level_tapbuf_size22_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_1_sram_inv[0:9]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size22 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_, chanx_right_in[5], chanx_right_in[19:20], chanx_right_in[34], chanx_left_in[10], chanx_left_in[25], chanx_left_in[35], chanx_left_in[40]}),
		.sram(mux_2level_tapbuf_size22_2_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_2_sram_inv[0:9]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size22 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_, chanx_right_in[6], chanx_right_in[21], chanx_right_in[23], chanx_right_in[36], chanx_left_in[9], chanx_left_in[24], chanx_left_in[31], chanx_left_in[38]}),
		.sram(mux_2level_tapbuf_size22_3_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_3_sram_inv[0:9]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size22 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_, chanx_right_in[0], chanx_right_in[3], chanx_right_in[14], chanx_right_in[29], chanx_left_in[1], chanx_left_in[7], chanx_left_in[16], chanx_left_in[30]}),
		.sram(mux_2level_tapbuf_size22_4_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_4_sram_inv[0:9]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size22 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[14], chany_top_in[29], chany_bottom_in[13], chany_bottom_in[28], chany_bottom_in[41], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size22_5_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_5_sram_inv[0:9]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size22 mux_left_track_9 (
		.in({chany_top_in[13], chany_top_in[28], chany_top_in[41], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[14], chany_bottom_in[29], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_}),
		.sram(mux_2level_tapbuf_size22_6_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_6_sram_inv[0:9]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size22 mux_left_track_17 (
		.in({chany_top_in[12], chany_top_in[26], chany_top_in[39], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[16], chany_bottom_in[30], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_}),
		.sram(mux_2level_tapbuf_size22_7_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_7_sram_inv[0:9]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size22 mux_left_track_33 (
		.in({chany_top_in[9], chany_top_in[24], chany_top_in[31], chany_top_in[38], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[18], chany_bottom_in[33], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_}),
		.sram(mux_2level_tapbuf_size22_8_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_8_sram_inv[0:9]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size22 mux_left_track_73 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[17], chany_top_in[32], chany_bottom_in[10], chany_bottom_in[25], chany_bottom_in[35], chany_bottom_in[40], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_}),
		.sram(mux_2level_tapbuf_size22_9_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size22_9_sram_inv[0:9]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size22_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_0_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_1_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_2_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_2_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_3_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_3_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size20_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_4_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_4_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_5_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_5_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_6_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_6_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_7_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_7_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_8_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_8_sram_inv[0:9]));

	mux_2level_tapbuf_size22_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size22_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size22_9_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size22_9_sram_inv[0:9]));

	mux_2level_tapbuf_size21 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[12], chanx_right_in[26], chanx_right_in[39], chanx_left_in[4], chanx_left_in[15], chanx_left_in[18], chanx_left_in[33]}),
		.sram(mux_2level_tapbuf_size21_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size21_0_sram_inv[0:9]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size21 mux_left_track_81 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[16], chany_top_in[30], chany_bottom_in[12], chany_bottom_in[26], chany_bottom_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_}),
		.sram(mux_2level_tapbuf_size21_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size21_1_sram_inv[0:9]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size21_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size23_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size21_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size21_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size21_0_sram_inv[0:9]));

	mux_2level_tapbuf_size21_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_9_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size21_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size21_1_sram_inv[0:9]));

	mux_2level_tapbuf_size20 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_, chanx_right_in[13], chanx_right_in[28], chanx_right_in[41], chanx_left_in[2], chanx_left_in[11], chanx_left_in[17], chanx_left_in[32]}),
		.sram(mux_2level_tapbuf_size20_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size20_0_sram_inv[0:9]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size20_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size21_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size20_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size20_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size20_0_sram_inv[0:9]));

	mux_2level_tapbuf_size6 mux_right_track_0 (
		.in({chany_top_in[13], chany_top_in[28], chany_top_in[41], chany_bottom_in[12], chany_bottom_in[26], chany_bottom_in[39]}),
		.sram(mux_2level_tapbuf_size6_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_0_sram_inv[0:5]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size6 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[26], chany_top_in[39], chany_bottom_in[13], chany_bottom_in[28], chany_bottom_in[41]}),
		.sram(mux_2level_tapbuf_size6_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_1_sram_inv[0:5]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size6_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size22_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_0_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[14], chany_top_in[29], chany_bottom_in[10], chany_bottom_in[25], chany_bottom_in[35], chany_bottom_in[40]}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size8 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[16], chany_top_in[30], chany_bottom_in[9], chany_bottom_in[24], chany_bottom_in[31], chany_bottom_in[38]}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size8 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[17], chany_top_in[32], chany_bottom_in[8], chany_bottom_in[22], chany_bottom_in[27], chany_bottom_in[37]}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size8 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[18], chany_top_in[33], chany_bottom_in[6], chany_bottom_in[21], chany_bottom_in[23], chany_bottom_in[36]}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size8 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19:20], chany_top_in[34], chany_bottom_in[5], chany_bottom_in[19:20], chany_bottom_in[34]}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size8 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[21], chany_top_in[23], chany_top_in[36], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[18], chany_bottom_in[33]}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size8 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[22], chany_top_in[27], chany_top_in[37], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[17], chany_bottom_in[32]}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size8 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[24], chany_top_in[31], chany_top_in[38], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[16], chany_bottom_in[30]}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size8 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[25], chany_top_in[35], chany_top_in[40], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[14], chany_bottom_in[29]}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size8 mux_bottom_track_9 (
		.in({chanx_right_in[10], chanx_right_in[25], chanx_right_in[35], chanx_right_in[40], chanx_left_in[2], chanx_left_in[11], chanx_left_in[17], chanx_left_in[32]}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size8 mux_bottom_track_17 (
		.in({chanx_right_in[9], chanx_right_in[24], chanx_right_in[31], chanx_right_in[38], chanx_left_in[4], chanx_left_in[15], chanx_left_in[18], chanx_left_in[33]}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size8 mux_bottom_track_25 (
		.in({chanx_right_in[8], chanx_right_in[22], chanx_right_in[27], chanx_right_in[37], chanx_left_in[5], chanx_left_in[19:20], chanx_left_in[34]}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size8 mux_bottom_track_33 (
		.in({chanx_right_in[6], chanx_right_in[21], chanx_right_in[23], chanx_right_in[36], chanx_left_in[6], chanx_left_in[21], chanx_left_in[23], chanx_left_in[36]}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size8 mux_bottom_track_41 (
		.in({chanx_right_in[5], chanx_right_in[19:20], chanx_right_in[34], chanx_left_in[8], chanx_left_in[22], chanx_left_in[27], chanx_left_in[37]}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size8 mux_bottom_track_49 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[18], chanx_right_in[33], chanx_left_in[9], chanx_left_in[24], chanx_left_in[31], chanx_left_in[38]}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size8 mux_bottom_track_57 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[17], chanx_right_in[32], chanx_left_in[10], chanx_left_in[25], chanx_left_in[35], chanx_left_in[40]}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size8_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size7 mux_bottom_track_1 (
		.in({chanx_right_in[12], chanx_right_in[26], chanx_right_in[39], chanx_left_in[1], chanx_left_in[7], chanx_left_in[16], chanx_left_in[30]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size7 mux_bottom_track_65 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[16], chanx_right_in[30], chanx_left_in[12], chanx_left_in[26], chanx_left_in[39]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size7 mux_bottom_track_73 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[14], chanx_right_in[29], chanx_left_in[13], chanx_left_in[28], chanx_left_in[41]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size7 mux_bottom_track_81 (
		.in({chanx_right_in[13], chanx_right_in[28], chanx_right_in[41], chanx_left_in[0], chanx_left_in[3], chanx_left_in[14], chanx_left_in[29]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

endmodule
// ----- END Verilog module for sb_4__3_ -----

//----- Default net type -----
`default_nettype wire



