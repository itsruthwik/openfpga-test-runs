//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug 20 23:36:48 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(pReset,
                prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:191] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:41] cbx_1__0__0_chanx_left_out;
wire [0:41] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:41] cbx_1__0__1_chanx_left_out;
wire [0:41] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:41] cbx_1__0__2_chanx_left_out;
wire [0:41] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:41] cbx_1__0__3_chanx_left_out;
wire [0:41] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:41] cbx_1__0__4_chanx_left_out;
wire [0:41] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:41] cbx_1__0__5_chanx_left_out;
wire [0:41] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:41] cbx_1__1__0_chanx_left_out;
wire [0:41] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:41] cbx_1__1__1_chanx_left_out;
wire [0:41] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__2_ccff_tail;
wire [0:41] cbx_1__1__2_chanx_left_out;
wire [0:41] cbx_1__1__2_chanx_right_out;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__3_ccff_tail;
wire [0:41] cbx_1__1__3_chanx_left_out;
wire [0:41] cbx_1__1__3_chanx_right_out;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__4_ccff_tail;
wire [0:41] cbx_1__1__4_chanx_left_out;
wire [0:41] cbx_1__1__4_chanx_right_out;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__5_ccff_tail;
wire [0:41] cbx_1__1__5_chanx_left_out;
wire [0:41] cbx_1__1__5_chanx_right_out;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:41] cbx_1__2__0_chanx_left_out;
wire [0:41] cbx_1__2__0_chanx_right_out;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:41] cbx_1__2__1_chanx_left_out;
wire [0:41] cbx_1__2__1_chanx_right_out;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__2_ccff_tail;
wire [0:41] cbx_1__2__2_chanx_left_out;
wire [0:41] cbx_1__2__2_chanx_right_out;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__3_ccff_tail;
wire [0:41] cbx_1__2__3_chanx_left_out;
wire [0:41] cbx_1__2__3_chanx_right_out;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__4_ccff_tail;
wire [0:41] cbx_1__2__4_chanx_left_out;
wire [0:41] cbx_1__2__4_chanx_right_out;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__2__5_ccff_tail;
wire [0:41] cbx_1__2__5_chanx_left_out;
wire [0:41] cbx_1__2__5_chanx_right_out;
wire [0:41] cbx_1__3__0_chanx_left_out;
wire [0:41] cbx_1__3__0_chanx_right_out;
wire [0:41] cbx_1__3__10_chanx_left_out;
wire [0:41] cbx_1__3__10_chanx_right_out;
wire [0:41] cbx_1__3__11_chanx_left_out;
wire [0:41] cbx_1__3__11_chanx_right_out;
wire [0:41] cbx_1__3__1_chanx_left_out;
wire [0:41] cbx_1__3__1_chanx_right_out;
wire [0:41] cbx_1__3__2_chanx_left_out;
wire [0:41] cbx_1__3__2_chanx_right_out;
wire [0:41] cbx_1__3__3_chanx_left_out;
wire [0:41] cbx_1__3__3_chanx_right_out;
wire [0:41] cbx_1__3__4_chanx_left_out;
wire [0:41] cbx_1__3__4_chanx_right_out;
wire [0:41] cbx_1__3__5_chanx_left_out;
wire [0:41] cbx_1__3__5_chanx_right_out;
wire [0:41] cbx_1__3__6_chanx_left_out;
wire [0:41] cbx_1__3__6_chanx_right_out;
wire [0:41] cbx_1__3__7_chanx_left_out;
wire [0:41] cbx_1__3__7_chanx_right_out;
wire [0:41] cbx_1__3__8_chanx_left_out;
wire [0:41] cbx_1__3__8_chanx_right_out;
wire [0:41] cbx_1__3__9_chanx_left_out;
wire [0:41] cbx_1__3__9_chanx_right_out;
wire [0:41] cbx_1__6__0_chanx_left_out;
wire [0:41] cbx_1__6__0_chanx_right_out;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__1_ccff_tail;
wire [0:41] cbx_1__6__1_chanx_left_out;
wire [0:41] cbx_1__6__1_chanx_right_out;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__2_ccff_tail;
wire [0:41] cbx_1__6__2_chanx_left_out;
wire [0:41] cbx_1__6__2_chanx_right_out;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__3_ccff_tail;
wire [0:41] cbx_1__6__3_chanx_left_out;
wire [0:41] cbx_1__6__3_chanx_right_out;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__3__0_ccff_tail;
wire [0:41] cbx_4__3__0_chanx_left_out;
wire [0:41] cbx_4__3__0_chanx_right_out;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_4__3__1_ccff_tail;
wire [0:41] cbx_4__3__1_chanx_left_out;
wire [0:41] cbx_4__3__1_chanx_right_out;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_4__3__2_ccff_tail;
wire [0:41] cbx_4__3__2_chanx_left_out;
wire [0:41] cbx_4__3__2_chanx_right_out;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_4__3__3_ccff_tail;
wire [0:41] cbx_4__3__3_chanx_left_out;
wire [0:41] cbx_4__3__3_chanx_right_out;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_4__4__0_ccff_tail;
wire [0:41] cbx_4__4__0_chanx_left_out;
wire [0:41] cbx_4__4__0_chanx_right_out;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_4__4__1_ccff_tail;
wire [0:41] cbx_4__4__1_chanx_left_out;
wire [0:41] cbx_4__4__1_chanx_right_out;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_4__6__0_ccff_tail;
wire [0:41] cbx_4__6__0_chanx_left_out;
wire [0:41] cbx_4__6__0_chanx_right_out;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_4__6__1_ccff_tail;
wire [0:41] cbx_4__6__1_chanx_left_out;
wire [0:41] cbx_4__6__1_chanx_right_out;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:41] cby_0__1__0_chany_bottom_out;
wire [0:41] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:41] cby_0__1__1_chany_bottom_out;
wire [0:41] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:41] cby_0__1__2_chany_bottom_out;
wire [0:41] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:41] cby_0__1__3_chany_bottom_out;
wire [0:41] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:41] cby_0__1__4_chany_bottom_out;
wire [0:41] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__2__0_ccff_tail;
wire [0:41] cby_0__2__0_chany_bottom_out;
wire [0:41] cby_0__2__0_chany_top_out;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:41] cby_1__1__0_chany_bottom_out;
wire [0:41] cby_1__1__0_chany_top_out;
wire [0:41] cby_1__1__10_chany_bottom_out;
wire [0:41] cby_1__1__10_chany_top_out;
wire [0:41] cby_1__1__11_chany_bottom_out;
wire [0:41] cby_1__1__11_chany_top_out;
wire [0:41] cby_1__1__12_chany_bottom_out;
wire [0:41] cby_1__1__12_chany_top_out;
wire [0:41] cby_1__1__13_chany_bottom_out;
wire [0:41] cby_1__1__13_chany_top_out;
wire [0:41] cby_1__1__14_chany_bottom_out;
wire [0:41] cby_1__1__14_chany_top_out;
wire [0:41] cby_1__1__15_chany_bottom_out;
wire [0:41] cby_1__1__15_chany_top_out;
wire [0:41] cby_1__1__16_chany_bottom_out;
wire [0:41] cby_1__1__16_chany_top_out;
wire [0:41] cby_1__1__17_chany_bottom_out;
wire [0:41] cby_1__1__17_chany_top_out;
wire [0:41] cby_1__1__18_chany_bottom_out;
wire [0:41] cby_1__1__18_chany_top_out;
wire [0:41] cby_1__1__1_chany_bottom_out;
wire [0:41] cby_1__1__1_chany_top_out;
wire [0:41] cby_1__1__2_chany_bottom_out;
wire [0:41] cby_1__1__2_chany_top_out;
wire [0:41] cby_1__1__3_chany_bottom_out;
wire [0:41] cby_1__1__3_chany_top_out;
wire [0:41] cby_1__1__4_chany_bottom_out;
wire [0:41] cby_1__1__4_chany_top_out;
wire [0:41] cby_1__1__5_chany_bottom_out;
wire [0:41] cby_1__1__5_chany_top_out;
wire [0:41] cby_1__1__6_chany_bottom_out;
wire [0:41] cby_1__1__6_chany_top_out;
wire [0:41] cby_1__1__7_chany_bottom_out;
wire [0:41] cby_1__1__7_chany_top_out;
wire [0:41] cby_1__1__8_chany_bottom_out;
wire [0:41] cby_1__1__8_chany_top_out;
wire [0:41] cby_1__1__9_chany_bottom_out;
wire [0:41] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__2__0_ccff_tail;
wire [0:41] cby_1__2__0_chany_bottom_out;
wire [0:41] cby_1__2__0_chany_top_out;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__1_ccff_tail;
wire [0:41] cby_1__2__1_chany_bottom_out;
wire [0:41] cby_1__2__1_chany_top_out;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__2_ccff_tail;
wire [0:41] cby_1__2__2_chany_bottom_out;
wire [0:41] cby_1__2__2_chany_top_out;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__3_ccff_tail;
wire [0:41] cby_1__2__3_chany_bottom_out;
wire [0:41] cby_1__2__3_chany_top_out;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__4_ccff_tail;
wire [0:41] cby_1__2__4_chany_bottom_out;
wire [0:41] cby_1__2__4_chany_top_out;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__4__0_ccff_tail;
wire [0:41] cby_3__4__0_chany_bottom_out;
wire [0:41] cby_3__4__0_chany_top_out;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_3__4__1_ccff_tail;
wire [0:41] cby_3__4__1_chany_bottom_out;
wire [0:41] cby_3__4__1_chany_top_out;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_3__4__2_ccff_tail;
wire [0:41] cby_3__4__2_chany_bottom_out;
wire [0:41] cby_3__4__2_chany_top_out;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_3__4__3_ccff_tail;
wire [0:41] cby_3__4__3_chany_bottom_out;
wire [0:41] cby_3__4__3_chany_top_out;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_4__4__0_ccff_tail;
wire [0:41] cby_4__4__0_chany_bottom_out;
wire [0:41] cby_4__4__0_chany_top_out;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_4__4__1_ccff_tail;
wire [0:41] cby_4__4__1_chany_bottom_out;
wire [0:41] cby_4__4__1_chany_top_out;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_6__1__0_ccff_tail;
wire [0:41] cby_6__1__0_chany_bottom_out;
wire [0:41] cby_6__1__0_chany_top_out;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_6__1__1_ccff_tail;
wire [0:41] cby_6__1__1_chany_bottom_out;
wire [0:41] cby_6__1__1_chany_top_out;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_6__1__2_ccff_tail;
wire [0:41] cby_6__1__2_chany_bottom_out;
wire [0:41] cby_6__1__2_chany_top_out;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_6__2__0_ccff_tail;
wire [0:41] cby_6__2__0_chany_bottom_out;
wire [0:41] cby_6__2__0_chany_top_out;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_6__4__0_ccff_tail;
wire [0:41] cby_6__4__0_chany_bottom_out;
wire [0:41] cby_6__4__0_chany_top_out;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__4__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_6__4__1_ccff_tail;
wire [0:41] cby_6__4__1_chany_bottom_out;
wire [0:41] cby_6__4__1_chany_top_out;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_6__4__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_2_ccff_tail;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_3_ccff_tail;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_4_ccff_tail;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_5_ccff_tail;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_2_ccff_tail;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_3_ccff_tail;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_4_ccff_tail;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_5_ccff_tail;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_2_ccff_tail;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_3_ccff_tail;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_4_ccff_tail;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_5_ccff_tail;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_4__4__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_4__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_6__4__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:41] sb_0__0__0_chanx_right_out;
wire [0:41] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:41] sb_0__1__0_chanx_right_out;
wire [0:41] sb_0__1__0_chany_bottom_out;
wire [0:41] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:41] sb_0__2__0_chanx_right_out;
wire [0:41] sb_0__2__0_chany_bottom_out;
wire [0:41] sb_0__2__0_chany_top_out;
wire [0:0] sb_0__3__0_ccff_tail;
wire [0:41] sb_0__3__0_chanx_right_out;
wire [0:41] sb_0__3__0_chany_bottom_out;
wire [0:41] sb_0__3__0_chany_top_out;
wire [0:0] sb_0__3__1_ccff_tail;
wire [0:41] sb_0__3__1_chanx_right_out;
wire [0:41] sb_0__3__1_chany_bottom_out;
wire [0:41] sb_0__3__1_chany_top_out;
wire [0:0] sb_0__3__2_ccff_tail;
wire [0:41] sb_0__3__2_chanx_right_out;
wire [0:41] sb_0__3__2_chany_bottom_out;
wire [0:41] sb_0__3__2_chany_top_out;
wire [0:0] sb_0__6__0_ccff_tail;
wire [0:41] sb_0__6__0_chanx_right_out;
wire [0:41] sb_0__6__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:41] sb_1__0__0_chanx_left_out;
wire [0:41] sb_1__0__0_chanx_right_out;
wire [0:41] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:41] sb_1__0__1_chanx_left_out;
wire [0:41] sb_1__0__1_chanx_right_out;
wire [0:41] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:41] sb_1__0__2_chanx_left_out;
wire [0:41] sb_1__0__2_chanx_right_out;
wire [0:41] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:41] sb_1__0__3_chanx_left_out;
wire [0:41] sb_1__0__3_chanx_right_out;
wire [0:41] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:41] sb_1__0__4_chanx_left_out;
wire [0:41] sb_1__0__4_chanx_right_out;
wire [0:41] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:41] sb_1__1__0_chanx_left_out;
wire [0:41] sb_1__1__0_chanx_right_out;
wire [0:41] sb_1__1__0_chany_bottom_out;
wire [0:41] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:41] sb_1__1__1_chanx_left_out;
wire [0:41] sb_1__1__1_chanx_right_out;
wire [0:41] sb_1__1__1_chany_bottom_out;
wire [0:41] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:41] sb_1__1__2_chanx_left_out;
wire [0:41] sb_1__1__2_chanx_right_out;
wire [0:41] sb_1__1__2_chany_bottom_out;
wire [0:41] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:41] sb_1__1__3_chanx_left_out;
wire [0:41] sb_1__1__3_chanx_right_out;
wire [0:41] sb_1__1__3_chany_bottom_out;
wire [0:41] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:41] sb_1__1__4_chanx_left_out;
wire [0:41] sb_1__1__4_chanx_right_out;
wire [0:41] sb_1__1__4_chany_bottom_out;
wire [0:41] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:41] sb_1__2__0_chanx_left_out;
wire [0:41] sb_1__2__0_chanx_right_out;
wire [0:41] sb_1__2__0_chany_bottom_out;
wire [0:41] sb_1__2__0_chany_top_out;
wire [0:0] sb_1__2__1_ccff_tail;
wire [0:41] sb_1__2__1_chanx_left_out;
wire [0:41] sb_1__2__1_chanx_right_out;
wire [0:41] sb_1__2__1_chany_bottom_out;
wire [0:41] sb_1__2__1_chany_top_out;
wire [0:0] sb_1__2__2_ccff_tail;
wire [0:41] sb_1__2__2_chanx_left_out;
wire [0:41] sb_1__2__2_chanx_right_out;
wire [0:41] sb_1__2__2_chany_bottom_out;
wire [0:41] sb_1__2__2_chany_top_out;
wire [0:0] sb_1__2__3_ccff_tail;
wire [0:41] sb_1__2__3_chanx_left_out;
wire [0:41] sb_1__2__3_chanx_right_out;
wire [0:41] sb_1__2__3_chany_bottom_out;
wire [0:41] sb_1__2__3_chany_top_out;
wire [0:0] sb_1__2__4_ccff_tail;
wire [0:41] sb_1__2__4_chanx_left_out;
wire [0:41] sb_1__2__4_chanx_right_out;
wire [0:41] sb_1__2__4_chany_bottom_out;
wire [0:41] sb_1__2__4_chany_top_out;
wire [0:0] sb_1__3__0_ccff_tail;
wire [0:41] sb_1__3__0_chanx_left_out;
wire [0:41] sb_1__3__0_chanx_right_out;
wire [0:41] sb_1__3__0_chany_bottom_out;
wire [0:41] sb_1__3__0_chany_top_out;
wire [0:0] sb_1__3__1_ccff_tail;
wire [0:41] sb_1__3__1_chanx_left_out;
wire [0:41] sb_1__3__1_chanx_right_out;
wire [0:41] sb_1__3__1_chany_bottom_out;
wire [0:41] sb_1__3__1_chany_top_out;
wire [0:0] sb_1__3__2_ccff_tail;
wire [0:41] sb_1__3__2_chanx_left_out;
wire [0:41] sb_1__3__2_chanx_right_out;
wire [0:41] sb_1__3__2_chany_bottom_out;
wire [0:41] sb_1__3__2_chany_top_out;
wire [0:0] sb_1__3__3_ccff_tail;
wire [0:41] sb_1__3__3_chanx_left_out;
wire [0:41] sb_1__3__3_chanx_right_out;
wire [0:41] sb_1__3__3_chany_bottom_out;
wire [0:41] sb_1__3__3_chany_top_out;
wire [0:0] sb_1__3__4_ccff_tail;
wire [0:41] sb_1__3__4_chanx_left_out;
wire [0:41] sb_1__3__4_chanx_right_out;
wire [0:41] sb_1__3__4_chany_bottom_out;
wire [0:41] sb_1__3__4_chany_top_out;
wire [0:0] sb_1__3__5_ccff_tail;
wire [0:41] sb_1__3__5_chanx_left_out;
wire [0:41] sb_1__3__5_chanx_right_out;
wire [0:41] sb_1__3__5_chany_bottom_out;
wire [0:41] sb_1__3__5_chany_top_out;
wire [0:0] sb_1__6__0_ccff_tail;
wire [0:41] sb_1__6__0_chanx_left_out;
wire [0:41] sb_1__6__0_chanx_right_out;
wire [0:41] sb_1__6__0_chany_bottom_out;
wire [0:0] sb_1__6__1_ccff_tail;
wire [0:41] sb_1__6__1_chanx_left_out;
wire [0:41] sb_1__6__1_chanx_right_out;
wire [0:41] sb_1__6__1_chany_bottom_out;
wire [0:0] sb_3__3__0_ccff_tail;
wire [0:41] sb_3__3__0_chanx_left_out;
wire [0:41] sb_3__3__0_chanx_right_out;
wire [0:41] sb_3__3__0_chany_bottom_out;
wire [0:41] sb_3__3__0_chany_top_out;
wire [0:0] sb_3__3__1_ccff_tail;
wire [0:41] sb_3__3__1_chanx_left_out;
wire [0:41] sb_3__3__1_chanx_right_out;
wire [0:41] sb_3__3__1_chany_bottom_out;
wire [0:41] sb_3__3__1_chany_top_out;
wire [0:0] sb_3__3__2_ccff_tail;
wire [0:41] sb_3__3__2_chanx_left_out;
wire [0:41] sb_3__3__2_chanx_right_out;
wire [0:41] sb_3__3__2_chany_bottom_out;
wire [0:41] sb_3__3__2_chany_top_out;
wire [0:0] sb_3__3__3_ccff_tail;
wire [0:41] sb_3__3__3_chanx_left_out;
wire [0:41] sb_3__3__3_chanx_right_out;
wire [0:41] sb_3__3__3_chany_bottom_out;
wire [0:41] sb_3__3__3_chany_top_out;
wire [0:0] sb_3__4__0_ccff_tail;
wire [0:41] sb_3__4__0_chanx_left_out;
wire [0:41] sb_3__4__0_chanx_right_out;
wire [0:41] sb_3__4__0_chany_bottom_out;
wire [0:41] sb_3__4__0_chany_top_out;
wire [0:0] sb_3__4__1_ccff_tail;
wire [0:41] sb_3__4__1_chanx_left_out;
wire [0:41] sb_3__4__1_chanx_right_out;
wire [0:41] sb_3__4__1_chany_bottom_out;
wire [0:41] sb_3__4__1_chany_top_out;
wire [0:0] sb_3__6__0_ccff_tail;
wire [0:41] sb_3__6__0_chanx_left_out;
wire [0:41] sb_3__6__0_chanx_right_out;
wire [0:41] sb_3__6__0_chany_bottom_out;
wire [0:0] sb_3__6__1_ccff_tail;
wire [0:41] sb_3__6__1_chanx_left_out;
wire [0:41] sb_3__6__1_chanx_right_out;
wire [0:41] sb_3__6__1_chany_bottom_out;
wire [0:0] sb_4__3__0_ccff_tail;
wire [0:41] sb_4__3__0_chanx_left_out;
wire [0:41] sb_4__3__0_chanx_right_out;
wire [0:41] sb_4__3__0_chany_bottom_out;
wire [0:41] sb_4__3__0_chany_top_out;
wire [0:0] sb_4__3__1_ccff_tail;
wire [0:41] sb_4__3__1_chanx_left_out;
wire [0:41] sb_4__3__1_chanx_right_out;
wire [0:41] sb_4__3__1_chany_bottom_out;
wire [0:41] sb_4__3__1_chany_top_out;
wire [0:0] sb_4__4__0_ccff_tail;
wire [0:41] sb_4__4__0_chanx_left_out;
wire [0:41] sb_4__4__0_chanx_right_out;
wire [0:41] sb_4__4__0_chany_bottom_out;
wire [0:41] sb_4__4__0_chany_top_out;
wire [0:0] sb_4__6__0_ccff_tail;
wire [0:41] sb_4__6__0_chanx_left_out;
wire [0:41] sb_4__6__0_chanx_right_out;
wire [0:41] sb_4__6__0_chany_bottom_out;
wire [0:0] sb_6__0__0_ccff_tail;
wire [0:41] sb_6__0__0_chanx_left_out;
wire [0:41] sb_6__0__0_chany_top_out;
wire [0:0] sb_6__1__0_ccff_tail;
wire [0:41] sb_6__1__0_chanx_left_out;
wire [0:41] sb_6__1__0_chany_bottom_out;
wire [0:41] sb_6__1__0_chany_top_out;
wire [0:0] sb_6__2__0_ccff_tail;
wire [0:41] sb_6__2__0_chanx_left_out;
wire [0:41] sb_6__2__0_chany_bottom_out;
wire [0:41] sb_6__2__0_chany_top_out;
wire [0:0] sb_6__3__0_ccff_tail;
wire [0:41] sb_6__3__0_chanx_left_out;
wire [0:41] sb_6__3__0_chany_bottom_out;
wire [0:41] sb_6__3__0_chany_top_out;
wire [0:0] sb_6__3__1_ccff_tail;
wire [0:41] sb_6__3__1_chanx_left_out;
wire [0:41] sb_6__3__1_chany_bottom_out;
wire [0:41] sb_6__3__1_chany_top_out;
wire [0:0] sb_6__4__0_ccff_tail;
wire [0:41] sb_6__4__0_chanx_left_out;
wire [0:41] sb_6__4__0_chany_bottom_out;
wire [0:41] sb_6__4__0_chany_top_out;
wire [0:0] sb_6__6__0_ccff_tail;
wire [0:41] sb_6__6__0_chanx_left_out;
wire [0:41] sb_6__6__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_top grid_io_top_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_top_5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_4_ccff_tail));

	grid_io_top grid_io_top_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_5_ccff_tail));

	grid_io_right grid_io_right_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right grid_io_right_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right grid_io_right_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_bottom grid_io_bottom_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[128:135]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_4_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[136:143]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_5_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[144:151]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[152:159]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__2__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[160:167]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[168:175]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[176:183]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[184:191]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__2__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__2__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__2__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__2__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_6__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_router grid_router_4__4_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_4__4__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	grid_router grid_router_4__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_4__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	grid_router grid_router_6__4_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__4__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	grid_router grid_router_6__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(ccff_head),
		.chany_top_out(sb_0__0__0_chany_top_out[0:41]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:41]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__2__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:41]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__2_ sb_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__2__0_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_0__2__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__2__0_chany_top_out[0:41]),
		.chanx_right_out(sb_0__2__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__2__0_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__2__0_ccff_tail));

	sb_0__3_ sb_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__3__0_chanx_left_out[0:41]),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__3__0_chany_top_out[0:41]),
		.chanx_right_out(sb_0__3__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__3__0_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__3__0_ccff_tail));

	sb_0__3_ sb_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__3__1_chanx_left_out[0:41]),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_0__3__1_chany_top_out[0:41]),
		.chanx_right_out(sb_0__3__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__3__1_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__3__1_ccff_tail));

	sb_0__3_ sb_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__3__2_chanx_left_out[0:41]),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_0__3__2_chany_top_out[0:41]),
		.chanx_right_out(sb_0__3__2_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__3__2_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__3__2_ccff_tail));

	sb_0__6_ sb_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__0_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__6__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_0__6__0_chany_bottom_out[0:41]),
		.ccff_tail(sb_0__6__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:41]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:41]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:41]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_bottom_5_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:41]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:41]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:41]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_bottom_4_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:41]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:41]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:41]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:41]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:41]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:41]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:41]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:41]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:41]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:41]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:41]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__1_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:41]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:41]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__2_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:41]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:41]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__3_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:41]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:41]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__4_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:41]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:41]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__2__1_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__2__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__0_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__2__0_chany_top_out[0:41]),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:41]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_1__2_ sb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__2__2_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__2__1_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__1_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__2__1_chany_top_out[0:41]),
		.chanx_right_out(sb_1__2__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__2__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__2__1_chanx_left_out[0:41]),
		.ccff_tail(sb_1__2__1_ccff_tail));

	sb_1__2_ sb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__2__3_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__2__2_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__2_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__2__2_chany_top_out[0:41]),
		.chanx_right_out(sb_1__2__2_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__2__2_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__2__2_chanx_left_out[0:41]),
		.ccff_tail(sb_1__2__2_ccff_tail));

	sb_1__2_ sb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__2__4_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__2__3_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__3_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__2__3_chany_top_out[0:41]),
		.chanx_right_out(sb_1__2__3_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__2__3_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__2__3_chanx_left_out[0:41]),
		.ccff_tail(sb_1__2__3_ccff_tail));

	sb_1__2_ sb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__2__5_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__2__4_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__4_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__2__4_chany_top_out[0:41]),
		.chanx_right_out(sb_1__2__4_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__2__4_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__2__4_chanx_left_out[0:41]),
		.ccff_tail(sb_1__2__4_ccff_tail));

	sb_1__3_ sb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__3_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__0_chanx_right_out[0:41]),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__3__0_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__0_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__0_ccff_tail));

	sb_1__3_ sb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__4_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__1_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__4_ccff_tail),
		.chany_top_out(sb_1__3__1_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__1_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__1_ccff_tail));

	sb_1__3_ sb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__5_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__2_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__1_ccff_tail),
		.chany_top_out(sb_1__3__2_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__2_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__2_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__2_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__2_ccff_tail));

	sb_1__3_ sb_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__6_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__3_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__0_ccff_tail),
		.chany_top_out(sb_1__3__3_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__3_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__3_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__3_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__3_ccff_tail));

	sb_1__3_ sb_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__7_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__4_chanx_right_out[0:41]),
		.ccff_head(cby_3__4__0_ccff_tail),
		.chany_top_out(sb_1__3__4_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__4_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__4_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__4_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__4_ccff_tail));

	sb_1__3_ sb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__8_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__5_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__2_ccff_tail),
		.chany_top_out(sb_1__3__5_chany_top_out[0:41]),
		.chanx_right_out(sb_1__3__5_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__3__5_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__3__5_chanx_left_out[0:41]),
		.ccff_tail(sb_1__3__5_ccff_tail));

	sb_1__6_ sb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__1_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__6__0_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__6__1_ccff_tail),
		.chanx_right_out(sb_1__6__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__6__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__6__0_chanx_left_out[0:41]),
		.ccff_tail(sb_1__6__0_ccff_tail));

	sb_1__6_ sb_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__2_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__6__1_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cby_3__4__1_ccff_tail),
		.chanx_right_out(sb_1__6__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_1__6__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_1__6__1_chanx_left_out[0:41]),
		.ccff_tail(sb_1__6__1_ccff_tail));

	sb_3__3_ sb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__4__0_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_4__3__0_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__6_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__3_ccff_tail),
		.chany_top_out(sb_3__3__0_chany_top_out[0:41]),
		.chanx_right_out(sb_3__3__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__3__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__3__0_chanx_left_out[0:41]),
		.ccff_tail(sb_3__3__0_ccff_tail));

	sb_3__3_ sb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__4__1_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_4__3__1_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__8_chanx_right_out[0:41]),
		.ccff_head(sb_1__3__5_ccff_tail),
		.chany_top_out(sb_3__3__1_chany_top_out[0:41]),
		.chanx_right_out(sb_3__3__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__3__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__3__1_chanx_left_out[0:41]),
		.ccff_tail(sb_3__3__1_ccff_tail));

	sb_3__3_ sb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__4__2_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_4__3__2_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__9_chanx_right_out[0:41]),
		.ccff_head(cbx_4__3__0_ccff_tail),
		.chany_top_out(sb_3__3__2_chany_top_out[0:41]),
		.chanx_right_out(sb_3__3__2_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__3__2_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__3__2_chanx_left_out[0:41]),
		.ccff_tail(sb_3__3__2_ccff_tail));

	sb_3__3_ sb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__4__3_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_4__3__3_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:41]),
		.chanx_left_in(cbx_1__3__11_chanx_right_out[0:41]),
		.ccff_head(cbx_4__3__1_ccff_tail),
		.chany_top_out(sb_3__3__3_chany_top_out[0:41]),
		.chanx_right_out(sb_3__3__3_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__3__3_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__3__3_chanx_left_out[0:41]),
		.ccff_tail(sb_3__3__3_ccff_tail));

	sb_3__4_ sb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_4__4__0_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_3__4__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_left_in(cbx_1__3__7_chanx_right_out[0:41]),
		.ccff_head(cby_4__4__0_ccff_tail),
		.chany_top_out(sb_3__4__0_chany_top_out[0:41]),
		.chanx_right_out(sb_3__4__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__4__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__4__0_chanx_left_out[0:41]),
		.ccff_tail(sb_3__4__0_ccff_tail));

	sb_3__4_ sb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_4__4__1_chanx_left_out[0:41]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_3__4__2_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_left_in(cbx_1__3__10_chanx_right_out[0:41]),
		.ccff_head(cby_6__4__0_ccff_tail),
		.chany_top_out(sb_3__4__1_chany_top_out[0:41]),
		.chanx_right_out(sb_3__4__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__4__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__4__1_chanx_left_out[0:41]),
		.ccff_tail(sb_3__4__1_ccff_tail));

	sb_3__6_ sb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_4__6__0_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_3__4__1_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_left_in(cbx_1__6__2_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cby_4__4__1_ccff_tail),
		.chanx_right_out(sb_3__6__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__6__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__6__0_chanx_left_out[0:41]),
		.ccff_tail(sb_3__6__0_ccff_tail));

	sb_3__6_ sb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_4__6__1_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_3__4__3_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_left_in(cbx_1__6__3_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cby_6__4__1_ccff_tail),
		.chanx_right_out(sb_3__6__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_3__6__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_3__6__1_chanx_left_out[0:41]),
		.ccff_tail(sb_3__6__1_ccff_tail));

	sb_4__3_ sb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__4__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_right_in(cbx_1__3__9_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:41]),
		.chanx_left_in(cbx_4__3__0_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.ccff_head(sb_3__3__0_ccff_tail),
		.chany_top_out(sb_4__3__0_chany_top_out[0:41]),
		.chanx_right_out(sb_4__3__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_4__3__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_4__3__0_chanx_left_out[0:41]),
		.ccff_tail(sb_4__3__0_ccff_tail));

	sb_4__3_ sb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__4__1_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_right_in(cbx_1__3__11_chanx_left_out[0:41]),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:41]),
		.chanx_left_in(cbx_4__3__1_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.ccff_head(sb_3__3__1_ccff_tail),
		.chany_top_out(sb_4__3__1_chany_top_out[0:41]),
		.chanx_right_out(sb_4__3__1_chanx_right_out[0:41]),
		.chany_bottom_out(sb_4__3__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_4__3__1_chanx_left_out[0:41]),
		.ccff_tail(sb_4__3__1_ccff_tail));

	sb_4__4_ sb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:41]),
		.chanx_right_in(cbx_1__3__10_chanx_left_out[0:41]),
		.chany_bottom_in(cby_4__4__0_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_4__4__0_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(cby_3__4__2_ccff_tail),
		.chany_top_out(sb_4__4__0_chany_top_out[0:41]),
		.chanx_right_out(sb_4__4__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_4__4__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_4__4__0_chanx_left_out[0:41]),
		.ccff_tail(sb_4__4__0_ccff_tail));

	sb_4__6_ sb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__3_chanx_left_out[0:41]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__4__1_chany_top_out[0:41]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_4__6__0_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(cby_3__4__3_ccff_tail),
		.chanx_right_out(sb_4__6__0_chanx_right_out[0:41]),
		.chany_bottom_out(sb_4__6__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_4__6__0_chanx_left_out[0:41]),
		.ccff_tail(sb_4__6__0_ccff_tail));

	sb_6__0_ sb_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__1__0_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.chany_top_out(sb_6__0__0_chany_top_out[0:41]),
		.chanx_left_out(sb_6__0__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__0__0_ccff_tail));

	sb_6__1_ sb_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__2__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_6__1__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_top_out(sb_6__1__0_chany_top_out[0:41]),
		.chany_bottom_out(sb_6__1__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__1__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__1__0_ccff_tail));

	sb_6__2_ sb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__1__1_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_6__2__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__2__5_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_6__1__0_ccff_tail),
		.chany_top_out(sb_6__2__0_chany_top_out[0:41]),
		.chany_bottom_out(sb_6__2__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__2__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__2__0_ccff_tail));

	sb_6__3_ sb_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__4__0_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_6__1__1_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_4__3__2_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.ccff_head(sb_3__3__2_ccff_tail),
		.chany_top_out(sb_6__3__0_chany_top_out[0:41]),
		.chany_bottom_out(sb_6__3__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__3__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__3__0_ccff_tail));

	sb_6__3_ sb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__4__1_chany_bottom_out[0:41]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_6__1__2_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_4__3__3_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.ccff_head(sb_3__3__3_ccff_tail),
		.chany_top_out(sb_6__3__1_chany_top_out[0:41]),
		.chany_bottom_out(sb_6__3__1_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__3__1_chanx_left_out[0:41]),
		.ccff_tail(sb_6__3__1_ccff_tail));

	sb_6__4_ sb_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__1__2_chany_bottom_out[0:41]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_6__4__0_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_4__4__1_chanx_right_out[0:41]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(cby_6__1__1_ccff_tail),
		.chany_top_out(sb_6__4__0_chany_top_out[0:41]),
		.chany_bottom_out(sb_6__4__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__4__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__4__0_ccff_tail));

	sb_6__6_ sb_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_6__4__1_chany_top_out[0:41]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_4__6__1_chanx_right_out[0:41]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(cby_6__1__2_ccff_tail),
		.chany_bottom_out(sb_6__6__0_chany_bottom_out[0:41]),
		.chanx_left_out(sb_6__6__0_chanx_left_out[0:41]),
		.ccff_tail(sb_6__6__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:41]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:41]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:41]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:41]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:41]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__0__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:41]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:41]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:41]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:41]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:41]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__1__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__2_ cbx_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:41]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__0_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__0_ccff_tail));

	cbx_1__2_ cbx_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__2__1_chanx_left_out[0:41]),
		.ccff_head(sb_1__2__1_ccff_tail),
		.chanx_left_out(cbx_1__2__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__1_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__1_ccff_tail));

	cbx_1__2_ cbx_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__2__2_chanx_left_out[0:41]),
		.ccff_head(sb_1__2__2_ccff_tail),
		.chanx_left_out(cbx_1__2__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__2_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__2_ccff_tail));

	cbx_1__2_ cbx_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__2__3_chanx_left_out[0:41]),
		.ccff_head(sb_1__2__3_ccff_tail),
		.chanx_left_out(cbx_1__2__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__3_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__3_ccff_tail));

	cbx_1__2_ cbx_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__3_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__2__4_chanx_left_out[0:41]),
		.ccff_head(sb_1__2__4_ccff_tail),
		.chanx_left_out(cbx_1__2__4_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__4_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__4_ccff_tail));

	cbx_1__2_ cbx_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__4_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__2__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__5_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__2__5_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__2__5_ccff_tail));

	cbx_1__3_ cbx_1__3_ (
		.chanx_left_in(sb_0__3__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__0_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__0_chanx_right_out[0:41]));

	cbx_1__3_ cbx_1__4_ (
		.chanx_left_in(sb_0__3__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__1_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__1_chanx_right_out[0:41]));

	cbx_1__3_ cbx_1__5_ (
		.chanx_left_in(sb_0__3__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__2_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__2_chanx_right_out[0:41]));

	cbx_1__3_ cbx_2__3_ (
		.chanx_left_in(sb_1__3__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__3_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__3_chanx_right_out[0:41]));

	cbx_1__3_ cbx_2__4_ (
		.chanx_left_in(sb_1__3__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__4_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__4_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__4_chanx_right_out[0:41]));

	cbx_1__3_ cbx_2__5_ (
		.chanx_left_in(sb_1__3__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__3__5_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__5_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__5_chanx_right_out[0:41]));

	cbx_1__3_ cbx_3__3_ (
		.chanx_left_in(sb_1__3__3_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__3__0_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__6_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__6_chanx_right_out[0:41]));

	cbx_1__3_ cbx_3__4_ (
		.chanx_left_in(sb_1__3__4_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__4__0_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__7_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__7_chanx_right_out[0:41]));

	cbx_1__3_ cbx_3__5_ (
		.chanx_left_in(sb_1__3__5_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__3__1_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__8_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__8_chanx_right_out[0:41]));

	cbx_1__3_ cbx_5__3_ (
		.chanx_left_in(sb_4__3__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__3__2_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__9_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__9_chanx_right_out[0:41]));

	cbx_1__3_ cbx_5__4_ (
		.chanx_left_in(sb_4__4__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__4__1_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__10_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__10_chanx_right_out[0:41]));

	cbx_1__3_ cbx_5__5_ (
		.chanx_left_in(sb_4__3__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__3__3_chanx_left_out[0:41]),
		.chanx_left_out(cbx_1__3__11_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__3__11_chanx_right_out[0:41]));

	cbx_1__6_ cbx_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__6__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__6__0_chanx_left_out[0:41]),
		.ccff_head(sb_1__6__0_ccff_tail),
		.chanx_left_out(cbx_1__6__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__6__0_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(ccff_tail));

	cbx_1__6_ cbx_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__6__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_1__6__1_chanx_left_out[0:41]),
		.ccff_head(sb_1__6__1_ccff_tail),
		.chanx_left_out(cbx_1__6__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__6__1_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__6__1_ccff_tail));

	cbx_1__6_ cbx_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__6__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__6__0_chanx_left_out[0:41]),
		.ccff_head(sb_3__6__0_ccff_tail),
		.chanx_left_out(cbx_1__6__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__6__2_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__6__2_ccff_tail));

	cbx_1__6_ cbx_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_4__6__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_3__6__1_chanx_left_out[0:41]),
		.ccff_head(sb_3__6__1_ccff_tail),
		.chanx_left_out(cbx_1__6__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_1__6__3_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__6__3_ccff_tail));

	cbx_4__3_ cbx_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__3__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_4__3__0_chanx_left_out[0:41]),
		.ccff_head(sb_4__3__0_ccff_tail),
		.chanx_left_out(cbx_4__3__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__3__0_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.ccff_tail(cbx_4__3__0_ccff_tail));

	cbx_4__3_ cbx_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__3__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_4__3__1_chanx_left_out[0:41]),
		.ccff_head(sb_4__3__1_ccff_tail),
		.chanx_left_out(cbx_4__3__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__3__1_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.ccff_tail(cbx_4__3__1_ccff_tail));

	cbx_4__3_ cbx_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__3__2_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__3__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__3__0_ccff_tail),
		.chanx_left_out(cbx_4__3__2_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__3__2_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.ccff_tail(cbx_4__3__2_ccff_tail));

	cbx_4__3_ cbx_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__3__3_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__3__1_chanx_left_out[0:41]),
		.ccff_head(sb_6__3__1_ccff_tail),
		.chanx_left_out(cbx_4__3__3_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__3__3_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_4__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.ccff_tail(cbx_4__3__3_ccff_tail));

	cbx_4__4_ cbx_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__4__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_4__4__0_chanx_left_out[0:41]),
		.ccff_head(sb_4__4__0_ccff_tail),
		.chanx_left_out(cbx_4__4__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__4__0_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_4__4__0_ccff_tail));

	cbx_4__4_ cbx_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__4__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__4__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__4__0_ccff_tail),
		.chanx_left_out(cbx_4__4__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__4__1_chanx_right_out[0:41]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_4__4__1_ccff_tail));

	cbx_4__6_ cbx_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__6__0_chanx_right_out[0:41]),
		.chanx_right_in(sb_4__6__0_chanx_left_out[0:41]),
		.ccff_head(sb_4__6__0_ccff_tail),
		.chanx_left_out(cbx_4__6__0_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__6__0_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_4__6__0_ccff_tail));

	cbx_4__6_ cbx_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__6__1_chanx_right_out[0:41]),
		.chanx_right_in(sb_6__6__0_chanx_left_out[0:41]),
		.ccff_head(sb_6__6__0_ccff_tail),
		.chanx_left_out(cbx_4__6__1_chanx_left_out[0:41]),
		.chanx_right_out(cbx_4__6__1_chanx_right_out[0:41]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_4__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_4__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_4__6__1_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:41]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:41]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__2__0_chany_top_out[0:41]),
		.chany_top_in(sb_0__3__0_chany_bottom_out[0:41]),
		.ccff_head(sb_0__3__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__0_chany_top_out[0:41]),
		.chany_top_in(sb_0__3__1_chany_bottom_out[0:41]),
		.ccff_head(sb_0__3__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__1_chany_top_out[0:41]),
		.chany_top_in(sb_0__3__2_chany_bottom_out[0:41]),
		.ccff_head(sb_0__3__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__2_chany_top_out[0:41]),
		.chany_top_in(sb_0__6__0_chany_bottom_out[0:41]),
		.ccff_head(sb_0__6__0_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__2_ cby_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:41]),
		.chany_top_in(sb_0__2__0_chany_bottom_out[0:41]),
		.ccff_head(sb_0__2__0_ccff_tail),
		.chany_bottom_out(cby_0__2__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_0__2__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__2__0_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:41]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:41]));

	cby_1__1_ cby_1__3_ (
		.chany_bottom_in(sb_1__2__0_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__0_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:41]));

	cby_1__1_ cby_1__4_ (
		.chany_bottom_in(sb_1__3__0_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__1_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:41]));

	cby_1__1_ cby_1__5_ (
		.chany_bottom_in(sb_1__3__1_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__2_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:41]));

	cby_1__1_ cby_1__6_ (
		.chany_bottom_in(sb_1__3__2_chany_top_out[0:41]),
		.chany_top_in(sb_1__6__0_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:41]));

	cby_1__1_ cby_2__1_ (
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:41]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:41]));

	cby_1__1_ cby_2__3_ (
		.chany_bottom_in(sb_1__2__1_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__3_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:41]));

	cby_1__1_ cby_2__4_ (
		.chany_bottom_in(sb_1__3__3_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__4_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:41]));

	cby_1__1_ cby_2__5_ (
		.chany_bottom_in(sb_1__3__4_chany_top_out[0:41]),
		.chany_top_in(sb_1__3__5_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:41]));

	cby_1__1_ cby_2__6_ (
		.chany_bottom_in(sb_1__3__5_chany_top_out[0:41]),
		.chany_top_in(sb_1__6__1_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:41]));

	cby_1__1_ cby_3__1_ (
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:41]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:41]));

	cby_1__1_ cby_3__3_ (
		.chany_bottom_in(sb_1__2__2_chany_top_out[0:41]),
		.chany_top_in(sb_3__3__0_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:41]));

	cby_1__1_ cby_3__5_ (
		.chany_bottom_in(sb_3__4__0_chany_top_out[0:41]),
		.chany_top_in(sb_3__3__1_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:41]));

	cby_1__1_ cby_4__1_ (
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:41]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:41]));

	cby_1__1_ cby_4__3_ (
		.chany_bottom_in(sb_1__2__3_chany_top_out[0:41]),
		.chany_top_in(sb_4__3__0_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:41]));

	cby_1__1_ cby_4__5_ (
		.chany_bottom_in(sb_4__4__0_chany_top_out[0:41]),
		.chany_top_in(sb_4__3__1_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:41]));

	cby_1__1_ cby_5__1_ (
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:41]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:41]));

	cby_1__1_ cby_5__3_ (
		.chany_bottom_in(sb_1__2__4_chany_top_out[0:41]),
		.chany_top_in(sb_3__3__2_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:41]));

	cby_1__1_ cby_5__5_ (
		.chany_bottom_in(sb_3__4__1_chany_top_out[0:41]),
		.chany_top_in(sb_3__3__3_chany_bottom_out[0:41]),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:41]));

	cby_1__2_ cby_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:41]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__0_ccff_tail),
		.chany_bottom_out(cby_1__2__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__2__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__2__0_ccff_tail));

	cby_1__2_ cby_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:41]),
		.chany_top_in(sb_1__2__1_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__1_ccff_tail),
		.chany_bottom_out(cby_1__2__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__2__1_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__2__1_ccff_tail));

	cby_1__2_ cby_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:41]),
		.chany_top_in(sb_1__2__2_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__2_ccff_tail),
		.chany_bottom_out(cby_1__2__2_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__2__2_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__2__2_ccff_tail));

	cby_1__2_ cby_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:41]),
		.chany_top_in(sb_1__2__3_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__3_ccff_tail),
		.chany_bottom_out(cby_1__2__3_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__2__3_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__2__3_ccff_tail));

	cby_1__2_ cby_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:41]),
		.chany_top_in(sb_1__2__4_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__4_ccff_tail),
		.chany_bottom_out(cby_1__2__4_chany_bottom_out[0:41]),
		.chany_top_out(cby_1__2__4_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__2__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__2__4_ccff_tail));

	cby_3__4_ cby_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__3__0_chany_top_out[0:41]),
		.chany_top_in(sb_3__4__0_chany_bottom_out[0:41]),
		.ccff_head(sb_3__4__0_ccff_tail),
		.chany_bottom_out(cby_3__4__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_3__4__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_3__4__0_ccff_tail));

	cby_3__4_ cby_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__3__1_chany_top_out[0:41]),
		.chany_top_in(sb_3__6__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__6__2_ccff_tail),
		.chany_bottom_out(cby_3__4__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_3__4__1_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_3__4__1_ccff_tail));

	cby_3__4_ cby_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__3__2_chany_top_out[0:41]),
		.chany_top_in(sb_3__4__1_chany_bottom_out[0:41]),
		.ccff_head(sb_3__4__1_ccff_tail),
		.chany_bottom_out(cby_3__4__2_chany_bottom_out[0:41]),
		.chany_top_out(cby_3__4__2_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_3__4__2_ccff_tail));

	cby_3__4_ cby_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__3__3_chany_top_out[0:41]),
		.chany_top_in(sb_3__6__1_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__6__3_ccff_tail),
		.chany_bottom_out(cby_3__4__3_chany_bottom_out[0:41]),
		.chany_top_out(cby_3__4__3_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_3__4__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_3__4__3_ccff_tail));

	cby_4__4_ cby_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__3__0_chany_top_out[0:41]),
		.chany_top_in(sb_4__4__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__4__0_ccff_tail),
		.chany_bottom_out(cby_4__4__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_4__4__0_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_4__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_4__4__0_ccff_tail));

	cby_4__4_ cby_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__3__1_chany_top_out[0:41]),
		.chany_top_in(sb_4__6__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__6__0_ccff_tail),
		.chany_bottom_out(cby_4__4__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_4__4__1_chany_top_out[0:41]),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_4__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_4__4__1_ccff_tail));

	cby_6__1_ cby_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__0__0_chany_top_out[0:41]),
		.chany_top_in(sb_6__1__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_6__1__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__1__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_6__1__0_ccff_tail));

	cby_6__1_ cby_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__2__0_chany_top_out[0:41]),
		.chany_top_in(sb_6__3__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__3__2_ccff_tail),
		.chany_bottom_out(cby_6__1__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__1__1_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_6__1__1_ccff_tail));

	cby_6__1_ cby_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__4__0_chany_top_out[0:41]),
		.chany_top_in(sb_6__3__1_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__3__3_ccff_tail),
		.chany_bottom_out(cby_6__1__2_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__1__2_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_6__1__2_ccff_tail));

	cby_6__2_ cby_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__1__0_chany_top_out[0:41]),
		.chany_top_in(sb_6__2__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_1__2__5_ccff_tail),
		.chany_bottom_out(cby_6__2__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__2__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_6__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_6__2__0_ccff_tail));

	cby_6__4_ cby_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__3__0_chany_top_out[0:41]),
		.chany_top_in(sb_6__4__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__4__1_ccff_tail),
		.chany_bottom_out(cby_6__4__0_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__4__0_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__4__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__4__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_6__4__0_ccff_tail));

	cby_6__4_ cby_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__3__1_chany_top_out[0:41]),
		.chany_top_in(sb_6__6__0_chany_bottom_out[0:41]),
		.ccff_head(cbx_4__6__1_ccff_tail),
		.chany_bottom_out(cby_6__4__1_chany_bottom_out[0:41]),
		.chany_top_out(cby_6__4__1_chany_top_out[0:41]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_6__4__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__4__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_6__4__1_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




