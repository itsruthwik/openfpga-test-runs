//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[2][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Sep 25 16:03:58 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_2__5_ -----
module sb_2__5_(pReset,
                prog_clk,
                chany_top_in,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_,
                chanx_left_in,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:228] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_;
//----- INPUT PORTS -----
input [0:228] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:228] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:228] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:228] chany_top_out;
//----- OUTPUT PORTS -----
output [0:228] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:228] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:228] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size10_0_sram;
wire [0:7] mux_2level_tapbuf_size10_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_1_sram;
wire [0:7] mux_2level_tapbuf_size10_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_2_sram;
wire [0:7] mux_2level_tapbuf_size10_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_3_sram;
wire [0:7] mux_2level_tapbuf_size10_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_4_sram;
wire [0:7] mux_2level_tapbuf_size10_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_5_sram;
wire [0:7] mux_2level_tapbuf_size10_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_6_sram;
wire [0:7] mux_2level_tapbuf_size10_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_7_sram;
wire [0:7] mux_2level_tapbuf_size10_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_8_sram;
wire [0:7] mux_2level_tapbuf_size10_8_sram_inv;
wire [0:0] mux_2level_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_8_ccff_tail;
wire [0:7] mux_2level_tapbuf_size11_0_sram;
wire [0:7] mux_2level_tapbuf_size11_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size11_mem_0_ccff_tail;
wire [0:7] mux_2level_tapbuf_size12_0_sram;
wire [0:7] mux_2level_tapbuf_size12_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size12_mem_0_ccff_tail;
wire [0:7] mux_2level_tapbuf_size13_0_sram;
wire [0:7] mux_2level_tapbuf_size13_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_10_sram;
wire [0:7] mux_2level_tapbuf_size13_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_11_sram;
wire [0:7] mux_2level_tapbuf_size13_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_12_sram;
wire [0:7] mux_2level_tapbuf_size13_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_1_sram;
wire [0:7] mux_2level_tapbuf_size13_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_2_sram;
wire [0:7] mux_2level_tapbuf_size13_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_3_sram;
wire [0:7] mux_2level_tapbuf_size13_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_4_sram;
wire [0:7] mux_2level_tapbuf_size13_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_5_sram;
wire [0:7] mux_2level_tapbuf_size13_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_6_sram;
wire [0:7] mux_2level_tapbuf_size13_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_7_sram;
wire [0:7] mux_2level_tapbuf_size13_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_8_sram;
wire [0:7] mux_2level_tapbuf_size13_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_9_sram;
wire [0:7] mux_2level_tapbuf_size13_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size14_0_sram;
wire [0:7] mux_2level_tapbuf_size14_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_10_sram;
wire [0:7] mux_2level_tapbuf_size14_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_11_sram;
wire [0:7] mux_2level_tapbuf_size14_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_12_sram;
wire [0:7] mux_2level_tapbuf_size14_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_13_sram;
wire [0:7] mux_2level_tapbuf_size14_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_14_sram;
wire [0:7] mux_2level_tapbuf_size14_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_15_sram;
wire [0:7] mux_2level_tapbuf_size14_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_16_sram;
wire [0:7] mux_2level_tapbuf_size14_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_17_sram;
wire [0:7] mux_2level_tapbuf_size14_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_18_sram;
wire [0:7] mux_2level_tapbuf_size14_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_19_sram;
wire [0:7] mux_2level_tapbuf_size14_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_1_sram;
wire [0:7] mux_2level_tapbuf_size14_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_20_sram;
wire [0:7] mux_2level_tapbuf_size14_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_21_sram;
wire [0:7] mux_2level_tapbuf_size14_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_22_sram;
wire [0:7] mux_2level_tapbuf_size14_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_23_sram;
wire [0:7] mux_2level_tapbuf_size14_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_24_sram;
wire [0:7] mux_2level_tapbuf_size14_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_25_sram;
wire [0:7] mux_2level_tapbuf_size14_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_26_sram;
wire [0:7] mux_2level_tapbuf_size14_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_27_sram;
wire [0:7] mux_2level_tapbuf_size14_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_28_sram;
wire [0:7] mux_2level_tapbuf_size14_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_29_sram;
wire [0:7] mux_2level_tapbuf_size14_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_2_sram;
wire [0:7] mux_2level_tapbuf_size14_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_30_sram;
wire [0:7] mux_2level_tapbuf_size14_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_31_sram;
wire [0:7] mux_2level_tapbuf_size14_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_32_sram;
wire [0:7] mux_2level_tapbuf_size14_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_33_sram;
wire [0:7] mux_2level_tapbuf_size14_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_34_sram;
wire [0:7] mux_2level_tapbuf_size14_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_35_sram;
wire [0:7] mux_2level_tapbuf_size14_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_36_sram;
wire [0:7] mux_2level_tapbuf_size14_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_37_sram;
wire [0:7] mux_2level_tapbuf_size14_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_38_sram;
wire [0:7] mux_2level_tapbuf_size14_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_39_sram;
wire [0:7] mux_2level_tapbuf_size14_39_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_3_sram;
wire [0:7] mux_2level_tapbuf_size14_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_40_sram;
wire [0:7] mux_2level_tapbuf_size14_40_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_41_sram;
wire [0:7] mux_2level_tapbuf_size14_41_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_42_sram;
wire [0:7] mux_2level_tapbuf_size14_42_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_4_sram;
wire [0:7] mux_2level_tapbuf_size14_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_5_sram;
wire [0:7] mux_2level_tapbuf_size14_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_6_sram;
wire [0:7] mux_2level_tapbuf_size14_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_7_sram;
wire [0:7] mux_2level_tapbuf_size14_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_8_sram;
wire [0:7] mux_2level_tapbuf_size14_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_9_sram;
wire [0:7] mux_2level_tapbuf_size14_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size14_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_9_ccff_tail;
wire [0:9] mux_2level_tapbuf_size17_0_sram;
wire [0:9] mux_2level_tapbuf_size17_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size17_1_sram;
wire [0:9] mux_2level_tapbuf_size17_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size17_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size17_mem_1_ccff_tail;
wire [0:9] mux_2level_tapbuf_size18_0_sram;
wire [0:9] mux_2level_tapbuf_size18_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_10_sram;
wire [0:9] mux_2level_tapbuf_size18_10_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_11_sram;
wire [0:9] mux_2level_tapbuf_size18_11_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_12_sram;
wire [0:9] mux_2level_tapbuf_size18_12_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_13_sram;
wire [0:9] mux_2level_tapbuf_size18_13_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_14_sram;
wire [0:9] mux_2level_tapbuf_size18_14_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_15_sram;
wire [0:9] mux_2level_tapbuf_size18_15_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_16_sram;
wire [0:9] mux_2level_tapbuf_size18_16_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_17_sram;
wire [0:9] mux_2level_tapbuf_size18_17_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_18_sram;
wire [0:9] mux_2level_tapbuf_size18_18_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_19_sram;
wire [0:9] mux_2level_tapbuf_size18_19_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_1_sram;
wire [0:9] mux_2level_tapbuf_size18_1_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_20_sram;
wire [0:9] mux_2level_tapbuf_size18_20_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_21_sram;
wire [0:9] mux_2level_tapbuf_size18_21_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_22_sram;
wire [0:9] mux_2level_tapbuf_size18_22_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_23_sram;
wire [0:9] mux_2level_tapbuf_size18_23_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_24_sram;
wire [0:9] mux_2level_tapbuf_size18_24_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_25_sram;
wire [0:9] mux_2level_tapbuf_size18_25_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_26_sram;
wire [0:9] mux_2level_tapbuf_size18_26_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_27_sram;
wire [0:9] mux_2level_tapbuf_size18_27_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_28_sram;
wire [0:9] mux_2level_tapbuf_size18_28_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_29_sram;
wire [0:9] mux_2level_tapbuf_size18_29_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_2_sram;
wire [0:9] mux_2level_tapbuf_size18_2_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_30_sram;
wire [0:9] mux_2level_tapbuf_size18_30_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_31_sram;
wire [0:9] mux_2level_tapbuf_size18_31_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_32_sram;
wire [0:9] mux_2level_tapbuf_size18_32_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_33_sram;
wire [0:9] mux_2level_tapbuf_size18_33_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_34_sram;
wire [0:9] mux_2level_tapbuf_size18_34_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_35_sram;
wire [0:9] mux_2level_tapbuf_size18_35_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_36_sram;
wire [0:9] mux_2level_tapbuf_size18_36_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_37_sram;
wire [0:9] mux_2level_tapbuf_size18_37_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_3_sram;
wire [0:9] mux_2level_tapbuf_size18_3_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_4_sram;
wire [0:9] mux_2level_tapbuf_size18_4_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_5_sram;
wire [0:9] mux_2level_tapbuf_size18_5_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_6_sram;
wire [0:9] mux_2level_tapbuf_size18_6_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_7_sram;
wire [0:9] mux_2level_tapbuf_size18_7_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_8_sram;
wire [0:9] mux_2level_tapbuf_size18_8_sram_inv;
wire [0:9] mux_2level_tapbuf_size18_9_sram;
wire [0:9] mux_2level_tapbuf_size18_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size18_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size18_mem_9_ccff_tail;
wire [0:9] mux_2level_tapbuf_size19_0_sram;
wire [0:9] mux_2level_tapbuf_size19_0_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_10_sram;
wire [0:9] mux_2level_tapbuf_size19_10_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_11_sram;
wire [0:9] mux_2level_tapbuf_size19_11_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_12_sram;
wire [0:9] mux_2level_tapbuf_size19_12_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_13_sram;
wire [0:9] mux_2level_tapbuf_size19_13_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_14_sram;
wire [0:9] mux_2level_tapbuf_size19_14_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_15_sram;
wire [0:9] mux_2level_tapbuf_size19_15_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_16_sram;
wire [0:9] mux_2level_tapbuf_size19_16_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_17_sram;
wire [0:9] mux_2level_tapbuf_size19_17_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_1_sram;
wire [0:9] mux_2level_tapbuf_size19_1_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_2_sram;
wire [0:9] mux_2level_tapbuf_size19_2_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_3_sram;
wire [0:9] mux_2level_tapbuf_size19_3_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_4_sram;
wire [0:9] mux_2level_tapbuf_size19_4_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_5_sram;
wire [0:9] mux_2level_tapbuf_size19_5_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_6_sram;
wire [0:9] mux_2level_tapbuf_size19_6_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_7_sram;
wire [0:9] mux_2level_tapbuf_size19_7_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_8_sram;
wire [0:9] mux_2level_tapbuf_size19_8_sram_inv;
wire [0:9] mux_2level_tapbuf_size19_9_sram;
wire [0:9] mux_2level_tapbuf_size19_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size19_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size19_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_16_sram;
wire [0:5] mux_2level_tapbuf_size8_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_17_sram;
wire [0:5] mux_2level_tapbuf_size8_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_18_sram;
wire [0:5] mux_2level_tapbuf_size8_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_19_sram;
wire [0:5] mux_2level_tapbuf_size8_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_20_sram;
wire [0:5] mux_2level_tapbuf_size8_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_21_sram;
wire [0:5] mux_2level_tapbuf_size8_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_22_sram;
wire [0:5] mux_2level_tapbuf_size8_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_23_sram;
wire [0:5] mux_2level_tapbuf_size8_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_24_sram;
wire [0:5] mux_2level_tapbuf_size8_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_25_sram;
wire [0:5] mux_2level_tapbuf_size8_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_26_sram;
wire [0:5] mux_2level_tapbuf_size8_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_27_sram;
wire [0:5] mux_2level_tapbuf_size8_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_28_sram;
wire [0:5] mux_2level_tapbuf_size8_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_29_sram;
wire [0:5] mux_2level_tapbuf_size8_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_30_sram;
wire [0:5] mux_2level_tapbuf_size8_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_31_sram;
wire [0:5] mux_2level_tapbuf_size8_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size9_0_sram;
wire [0:7] mux_2level_tapbuf_size9_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_10_sram;
wire [0:7] mux_2level_tapbuf_size9_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_11_sram;
wire [0:7] mux_2level_tapbuf_size9_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_12_sram;
wire [0:7] mux_2level_tapbuf_size9_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_13_sram;
wire [0:7] mux_2level_tapbuf_size9_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_14_sram;
wire [0:7] mux_2level_tapbuf_size9_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_15_sram;
wire [0:7] mux_2level_tapbuf_size9_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_16_sram;
wire [0:7] mux_2level_tapbuf_size9_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_17_sram;
wire [0:7] mux_2level_tapbuf_size9_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_18_sram;
wire [0:7] mux_2level_tapbuf_size9_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_19_sram;
wire [0:7] mux_2level_tapbuf_size9_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_1_sram;
wire [0:7] mux_2level_tapbuf_size9_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_20_sram;
wire [0:7] mux_2level_tapbuf_size9_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_21_sram;
wire [0:7] mux_2level_tapbuf_size9_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_22_sram;
wire [0:7] mux_2level_tapbuf_size9_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_23_sram;
wire [0:7] mux_2level_tapbuf_size9_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_24_sram;
wire [0:7] mux_2level_tapbuf_size9_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_25_sram;
wire [0:7] mux_2level_tapbuf_size9_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_26_sram;
wire [0:7] mux_2level_tapbuf_size9_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_27_sram;
wire [0:7] mux_2level_tapbuf_size9_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_28_sram;
wire [0:7] mux_2level_tapbuf_size9_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_29_sram;
wire [0:7] mux_2level_tapbuf_size9_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_2_sram;
wire [0:7] mux_2level_tapbuf_size9_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_30_sram;
wire [0:7] mux_2level_tapbuf_size9_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_31_sram;
wire [0:7] mux_2level_tapbuf_size9_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_32_sram;
wire [0:7] mux_2level_tapbuf_size9_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_33_sram;
wire [0:7] mux_2level_tapbuf_size9_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_34_sram;
wire [0:7] mux_2level_tapbuf_size9_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_35_sram;
wire [0:7] mux_2level_tapbuf_size9_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_36_sram;
wire [0:7] mux_2level_tapbuf_size9_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_37_sram;
wire [0:7] mux_2level_tapbuf_size9_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_38_sram;
wire [0:7] mux_2level_tapbuf_size9_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_39_sram;
wire [0:7] mux_2level_tapbuf_size9_39_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_3_sram;
wire [0:7] mux_2level_tapbuf_size9_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_40_sram;
wire [0:7] mux_2level_tapbuf_size9_40_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_41_sram;
wire [0:7] mux_2level_tapbuf_size9_41_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_42_sram;
wire [0:7] mux_2level_tapbuf_size9_42_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_43_sram;
wire [0:7] mux_2level_tapbuf_size9_43_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_44_sram;
wire [0:7] mux_2level_tapbuf_size9_44_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_45_sram;
wire [0:7] mux_2level_tapbuf_size9_45_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_46_sram;
wire [0:7] mux_2level_tapbuf_size9_46_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_47_sram;
wire [0:7] mux_2level_tapbuf_size9_47_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_48_sram;
wire [0:7] mux_2level_tapbuf_size9_48_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_49_sram;
wire [0:7] mux_2level_tapbuf_size9_49_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_4_sram;
wire [0:7] mux_2level_tapbuf_size9_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_50_sram;
wire [0:7] mux_2level_tapbuf_size9_50_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_51_sram;
wire [0:7] mux_2level_tapbuf_size9_51_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_52_sram;
wire [0:7] mux_2level_tapbuf_size9_52_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_53_sram;
wire [0:7] mux_2level_tapbuf_size9_53_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_54_sram;
wire [0:7] mux_2level_tapbuf_size9_54_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_55_sram;
wire [0:7] mux_2level_tapbuf_size9_55_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_56_sram;
wire [0:7] mux_2level_tapbuf_size9_56_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_57_sram;
wire [0:7] mux_2level_tapbuf_size9_57_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_58_sram;
wire [0:7] mux_2level_tapbuf_size9_58_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_59_sram;
wire [0:7] mux_2level_tapbuf_size9_59_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_5_sram;
wire [0:7] mux_2level_tapbuf_size9_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_60_sram;
wire [0:7] mux_2level_tapbuf_size9_60_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_61_sram;
wire [0:7] mux_2level_tapbuf_size9_61_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_62_sram;
wire [0:7] mux_2level_tapbuf_size9_62_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_63_sram;
wire [0:7] mux_2level_tapbuf_size9_63_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_64_sram;
wire [0:7] mux_2level_tapbuf_size9_64_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_65_sram;
wire [0:7] mux_2level_tapbuf_size9_65_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_66_sram;
wire [0:7] mux_2level_tapbuf_size9_66_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_67_sram;
wire [0:7] mux_2level_tapbuf_size9_67_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_68_sram;
wire [0:7] mux_2level_tapbuf_size9_68_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_69_sram;
wire [0:7] mux_2level_tapbuf_size9_69_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_6_sram;
wire [0:7] mux_2level_tapbuf_size9_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_70_sram;
wire [0:7] mux_2level_tapbuf_size9_70_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_71_sram;
wire [0:7] mux_2level_tapbuf_size9_71_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_72_sram;
wire [0:7] mux_2level_tapbuf_size9_72_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_73_sram;
wire [0:7] mux_2level_tapbuf_size9_73_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_74_sram;
wire [0:7] mux_2level_tapbuf_size9_74_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_7_sram;
wire [0:7] mux_2level_tapbuf_size9_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_8_sram;
wire [0:7] mux_2level_tapbuf_size9_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_9_sram;
wire [0:7] mux_2level_tapbuf_size9_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[193] = chany_top_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[194] = chany_top_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[195] = chany_top_in[194];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[197] = chany_top_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[198] = chany_top_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[199] = chany_top_in[198];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[201] = chany_top_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[202] = chany_top_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[203] = chany_top_in[202];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[205] = chany_top_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[206] = chany_top_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[207] = chany_top_in[206];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[209] = chany_top_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[210] = chany_top_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[211] = chany_top_in[210];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[213] = chany_top_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[214] = chany_top_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[215] = chany_top_in[214];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[217] = chany_top_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[218] = chany_top_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[219] = chany_top_in[218];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[221] = chany_top_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[222] = chany_top_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[223] = chany_top_in[222];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[225] = chany_top_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[226] = chany_top_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[227] = chany_top_in[226];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[177] = chanx_right_in[176];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[178] = chanx_right_in[177];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[179] = chanx_right_in[178];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[181] = chanx_right_in[180];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[182] = chanx_right_in[181];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[183] = chanx_right_in[182];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[185] = chanx_right_in[184];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[186] = chanx_right_in[185];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[187] = chanx_right_in[186];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[189] = chanx_right_in[188];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[190] = chanx_right_in[189];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[191] = chanx_right_in[190];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[193] = chanx_right_in[192];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[194] = chanx_right_in[193];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[195] = chanx_right_in[194];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[197] = chanx_right_in[196];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[198] = chanx_right_in[197];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[199] = chanx_right_in[198];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[201] = chanx_right_in[200];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[202] = chanx_right_in[201];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[203] = chanx_right_in[202];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[205] = chanx_right_in[204];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[206] = chanx_right_in[205];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[207] = chanx_right_in[206];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[209] = chanx_right_in[208];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[210] = chanx_right_in[209];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[211] = chanx_right_in[210];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[213] = chanx_right_in[212];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[214] = chanx_right_in[213];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[215] = chanx_right_in[214];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[217] = chanx_right_in[216];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[218] = chanx_right_in[217];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[219] = chanx_right_in[218];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[221] = chanx_right_in[220];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[222] = chanx_right_in[221];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[223] = chanx_right_in[222];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[225] = chanx_right_in[224];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[226] = chanx_right_in[225];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[227] = chanx_right_in[226];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 713 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 714 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 717 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 718 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 721 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 722 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 725 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 726 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 729 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 730 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 733 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 734 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 737 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 738 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 741 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 742 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 745 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 746 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 749 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 750 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 753 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 754 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 757 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 758 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 761 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 762 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 765 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 766 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 769 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 770 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 773 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 774 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 777 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 778 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 781 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 782 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[193] = chany_bottom_in[192];
// ----- Local connection due to Wire 785 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[194] = chany_bottom_in[193];
// ----- Local connection due to Wire 786 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[195] = chany_bottom_in[194];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chany_bottom_in[196];
// ----- Local connection due to Wire 789 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[198] = chany_bottom_in[197];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[199] = chany_bottom_in[198];
// ----- Local connection due to Wire 792 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[201] = chany_bottom_in[200];
// ----- Local connection due to Wire 793 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[202] = chany_bottom_in[201];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[203] = chany_bottom_in[202];
// ----- Local connection due to Wire 796 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[205] = chany_bottom_in[204];
// ----- Local connection due to Wire 797 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chany_bottom_in[205];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[207] = chany_bottom_in[206];
// ----- Local connection due to Wire 800 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[209] = chany_bottom_in[208];
// ----- Local connection due to Wire 801 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[210] = chany_bottom_in[209];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[211] = chany_bottom_in[210];
// ----- Local connection due to Wire 804 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[213] = chany_bottom_in[212];
// ----- Local connection due to Wire 805 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[214] = chany_bottom_in[213];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chany_bottom_in[214];
// ----- Local connection due to Wire 808 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[217] = chany_bottom_in[216];
// ----- Local connection due to Wire 809 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[218] = chany_bottom_in[217];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[219] = chany_bottom_in[218];
// ----- Local connection due to Wire 812 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[221] = chany_bottom_in[220];
// ----- Local connection due to Wire 813 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[222] = chany_bottom_in[221];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[223] = chany_bottom_in[222];
// ----- Local connection due to Wire 816 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[225] = chany_bottom_in[224];
// ----- Local connection due to Wire 817 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[226] = chany_bottom_in[225];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[227] = chany_bottom_in[226];
// ----- Local connection due to Wire 831 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 832 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 833 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 835 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 836 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 837 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 839 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 840 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 841 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 843 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 844 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 845 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 847 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 848 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 849 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 851 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 852 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 853 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 855 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 856 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 857 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 859 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 860 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 861 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 863 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 864 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 865 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 867 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 868 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 869 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 871 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 872 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 873 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 875 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 876 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 877 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 879 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 880 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 881 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 883 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 884 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 885 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 887 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 888 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 889 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 891 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 892 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 893 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 895 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 896 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 897 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 899 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 900 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 901 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 903 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 904 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 905 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 907 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 908 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 909 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 911 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 912 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 913 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 915 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 916 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 917 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 919 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 920 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 921 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 923 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 924 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 925 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 927 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 928 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 929 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 931 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 932 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 933 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 935 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 936 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 937 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 939 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 940 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 941 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 943 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 944 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 945 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 947 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 948 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 949 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 951 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 952 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 953 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 955 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 956 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 957 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 959 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 960 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 961 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 963 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 964 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 965 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 967 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 968 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 969 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 971 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 972 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 973 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 975 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 976 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 977 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 979 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 980 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 981 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 983 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 984 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 985 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 987 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 988 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 989 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 991 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 992 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 993 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 995 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 996 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 997 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 999 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 1000 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 1001 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 1003 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 1004 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 1005 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- Local connection due to Wire 1007 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[177] = chanx_left_in[176];
// ----- Local connection due to Wire 1008 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[178] = chanx_left_in[177];
// ----- Local connection due to Wire 1009 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[179] = chanx_left_in[178];
// ----- Local connection due to Wire 1011 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[181] = chanx_left_in[180];
// ----- Local connection due to Wire 1012 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[182] = chanx_left_in[181];
// ----- Local connection due to Wire 1013 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[183] = chanx_left_in[182];
// ----- Local connection due to Wire 1015 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[185] = chanx_left_in[184];
// ----- Local connection due to Wire 1016 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[186] = chanx_left_in[185];
// ----- Local connection due to Wire 1017 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[187] = chanx_left_in[186];
// ----- Local connection due to Wire 1019 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[189] = chanx_left_in[188];
// ----- Local connection due to Wire 1020 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[190] = chanx_left_in[189];
// ----- Local connection due to Wire 1021 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[191] = chanx_left_in[190];
// ----- Local connection due to Wire 1023 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[193] = chanx_left_in[192];
// ----- Local connection due to Wire 1024 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[194] = chanx_left_in[193];
// ----- Local connection due to Wire 1025 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[195] = chanx_left_in[194];
// ----- Local connection due to Wire 1027 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[197] = chanx_left_in[196];
// ----- Local connection due to Wire 1028 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[198] = chanx_left_in[197];
// ----- Local connection due to Wire 1029 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[199] = chanx_left_in[198];
// ----- Local connection due to Wire 1031 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[201] = chanx_left_in[200];
// ----- Local connection due to Wire 1032 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[202] = chanx_left_in[201];
// ----- Local connection due to Wire 1033 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[203] = chanx_left_in[202];
// ----- Local connection due to Wire 1035 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[205] = chanx_left_in[204];
// ----- Local connection due to Wire 1036 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[206] = chanx_left_in[205];
// ----- Local connection due to Wire 1037 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[207] = chanx_left_in[206];
// ----- Local connection due to Wire 1039 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[209] = chanx_left_in[208];
// ----- Local connection due to Wire 1040 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[210] = chanx_left_in[209];
// ----- Local connection due to Wire 1041 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[211] = chanx_left_in[210];
// ----- Local connection due to Wire 1043 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[213] = chanx_left_in[212];
// ----- Local connection due to Wire 1044 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[214] = chanx_left_in[213];
// ----- Local connection due to Wire 1045 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[215] = chanx_left_in[214];
// ----- Local connection due to Wire 1047 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[217] = chanx_left_in[216];
// ----- Local connection due to Wire 1048 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[218] = chanx_left_in[217];
// ----- Local connection due to Wire 1049 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[219] = chanx_left_in[218];
// ----- Local connection due to Wire 1051 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[221] = chanx_left_in[220];
// ----- Local connection due to Wire 1052 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[222] = chanx_left_in[221];
// ----- Local connection due to Wire 1053 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[223] = chanx_left_in[222];
// ----- Local connection due to Wire 1055 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[225] = chanx_left_in[224];
// ----- Local connection due to Wire 1056 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[226] = chanx_left_in[225];
// ----- Local connection due to Wire 1057 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[227] = chanx_left_in[226];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size19 mux_top_track_0 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[78], chanx_right_in[156], chanx_left_in[0], chanx_left_in[3], chanx_left_in[77], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size19_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_0_sram_inv[0:9]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size19 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[6], chanx_right_in[23], chanx_right_in[84], chanx_right_in[161], chanx_left_in[72], chanx_left_in[149], chanx_left_in[219], chanx_left_in[226]}),
		.sram(mux_2level_tapbuf_size19_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_1_sram_inv[0:9]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size19 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[85], chanx_right_in[162], chanx_left_in[70], chanx_left_in[148], chanx_left_in[215], chanx_left_in[225]}),
		.sram(mux_2level_tapbuf_size19_2_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_2_sram_inv[0:9]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size19 mux_top_track_72 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[13], chanx_right_in[43], chanx_right_in[90], chanx_right_in[168], chanx_left_in[65], chanx_left_in[142], chanx_left_in[199], chanx_left_in[220]}),
		.sram(mux_2level_tapbuf_size19_3_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_3_sram_inv[0:9]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size19 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[14], chanx_right_in[47], chanx_right_in[92], chanx_right_in[169], chanx_left_in[64], chanx_left_in[141], chanx_left_in[195], chanx_left_in[218]}),
		.sram(mux_2level_tapbuf_size19_4_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_4_sram_inv[0:9]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size19 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[16], chanx_right_in[51], chanx_right_in[93], chanx_right_in[170], chanx_left_in[62], chanx_left_in[140], chanx_left_in[191], chanx_left_in[217]}),
		.sram(mux_2level_tapbuf_size19_5_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_5_sram_inv[0:9]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size19 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[17], chanx_right_in[55], chanx_right_in[94], chanx_right_in[172], chanx_left_in[61], chanx_left_in[138], chanx_left_in[187], chanx_left_in[216]}),
		.sram(mux_2level_tapbuf_size19_6_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_6_sram_inv[0:9]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size19 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[18], chanx_right_in[59], chanx_right_in[96], chanx_right_in[173], chanx_left_in[60], chanx_left_in[137], chanx_left_in[183], chanx_left_in[214]}),
		.sram(mux_2level_tapbuf_size19_7_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_7_sram_inv[0:9]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size19 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[20], chanx_right_in[63], chanx_right_in[97], chanx_right_in[174], chanx_left_in[58], chanx_left_in[136], chanx_left_in[179], chanx_left_in[213]}),
		.sram(mux_2level_tapbuf_size19_8_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_8_sram_inv[0:9]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size19 mux_top_track_144 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[25], chanx_right_in[79], chanx_right_in[102], chanx_right_in[180], chanx_left_in[53], chanx_left_in[130], chanx_left_in[163], chanx_left_in[208]}),
		.sram(mux_2level_tapbuf_size19_9_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_9_sram_inv[0:9]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size19 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[26], chanx_right_in[83], chanx_right_in[104], chanx_right_in[181], chanx_left_in[52], chanx_left_in[129], chanx_left_in[159], chanx_left_in[206]}),
		.sram(mux_2level_tapbuf_size19_10_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_10_sram_inv[0:9]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size19 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[28], chanx_right_in[87], chanx_right_in[105], chanx_right_in[182], chanx_left_in[50], chanx_left_in[128], chanx_left_in[155], chanx_left_in[205]}),
		.sram(mux_2level_tapbuf_size19_11_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_11_sram_inv[0:9]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size19 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[29], chanx_right_in[91], chanx_right_in[106], chanx_right_in[184], chanx_left_in[49], chanx_left_in[126], chanx_left_in[151], chanx_left_in[204]}),
		.sram(mux_2level_tapbuf_size19_12_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_12_sram_inv[0:9]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size19 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[30], chanx_right_in[95], chanx_right_in[108], chanx_right_in[185], chanx_left_in[48], chanx_left_in[125], chanx_left_in[147], chanx_left_in[202]}),
		.sram(mux_2level_tapbuf_size19_13_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_13_sram_inv[0:9]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size19 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[32], chanx_right_in[99], chanx_right_in[109], chanx_right_in[186], chanx_left_in[46], chanx_left_in[124], chanx_left_in[143], chanx_left_in[201]}),
		.sram(mux_2level_tapbuf_size19_14_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_14_sram_inv[0:9]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size19 mux_top_track_216 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[37], chanx_right_in[114:115], chanx_right_in[192], chanx_left_in[41], chanx_left_in[118], chanx_left_in[127], chanx_left_in[196]}),
		.sram(mux_2level_tapbuf_size19_15_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_15_sram_inv[0:9]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size19 mux_top_track_288 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[49], chanx_right_in[126], chanx_right_in[151], chanx_right_in[204], chanx_left_in[29], chanx_left_in[91], chanx_left_in[106], chanx_left_in[184]}),
		.sram(mux_2level_tapbuf_size19_16_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_16_sram_inv[0:9]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size19 mux_top_track_360 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[61], chanx_right_in[138], chanx_right_in[187], chanx_right_in[216], chanx_left_in[17], chanx_left_in[55], chanx_left_in[94], chanx_left_in[172]}),
		.sram(mux_2level_tapbuf_size19_17_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size19_17_sram_inv[0:9]),
		.out(chany_top_out[180]));

	mux_2level_tapbuf_size19_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size19_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_0_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_1_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_2_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_2_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_3_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_3_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_4_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_4_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_5_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_5_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_6_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_6_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_7_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_7_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_8_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_8_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_9_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_9_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_10_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_10_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_11_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_11_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_12_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_12_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_13_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_13_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_14_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_14_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_15_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_15_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_16_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_16_sram_inv[0:9]));

	mux_2level_tapbuf_size19_mem mem_top_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size19_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size19_17_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size19_17_sram_inv[0:9]));

	mux_2level_tapbuf_size18 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[80], chanx_right_in[157], chanx_left_in[76], chanx_left_in[153], chanx_left_in[228]}),
		.sram(mux_2level_tapbuf_size18_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_0_sram_inv[0:9]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size18 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[4], chanx_right_in[15], chanx_right_in[81], chanx_right_in[158], chanx_left_in[74], chanx_left_in[152], chanx_left_in[227]}),
		.sram(mux_2level_tapbuf_size18_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_1_sram_inv[0:9]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size18 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[5], chanx_right_in[19], chanx_right_in[82], chanx_right_in[160], chanx_left_in[73], chanx_left_in[150], chanx_left_in[223]}),
		.sram(mux_2level_tapbuf_size18_2_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_2_sram_inv[0:9]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size18 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[9], chanx_right_in[31], chanx_right_in[86], chanx_right_in[164], chanx_left_in[69], chanx_left_in[146], chanx_left_in[211], chanx_left_in[224]}),
		.sram(mux_2level_tapbuf_size18_3_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_3_sram_inv[0:9]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size18 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[10], chanx_right_in[35], chanx_right_in[88], chanx_right_in[165], chanx_left_in[68], chanx_left_in[145], chanx_left_in[207], chanx_left_in[222]}),
		.sram(mux_2level_tapbuf_size18_4_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_4_sram_inv[0:9]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size18 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[12], chanx_right_in[39], chanx_right_in[89], chanx_right_in[166], chanx_left_in[66], chanx_left_in[144], chanx_left_in[203], chanx_left_in[221]}),
		.sram(mux_2level_tapbuf_size18_5_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_5_sram_inv[0:9]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size18 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[21], chanx_right_in[67], chanx_right_in[98], chanx_right_in[176], chanx_left_in[57], chanx_left_in[134], chanx_left_in[175], chanx_left_in[212]}),
		.sram(mux_2level_tapbuf_size18_6_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_6_sram_inv[0:9]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size18 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[22], chanx_right_in[71], chanx_right_in[100], chanx_right_in[177], chanx_left_in[56], chanx_left_in[133], chanx_left_in[171], chanx_left_in[210]}),
		.sram(mux_2level_tapbuf_size18_7_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_7_sram_inv[0:9]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size18 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[24], chanx_right_in[75], chanx_right_in[101], chanx_right_in[178], chanx_left_in[54], chanx_left_in[132], chanx_left_in[167], chanx_left_in[209]}),
		.sram(mux_2level_tapbuf_size18_8_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_8_sram_inv[0:9]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size18 mux_top_track_192 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[33], chanx_right_in[103], chanx_right_in[110], chanx_right_in[188], chanx_left_in[45], chanx_left_in[122], chanx_left_in[139], chanx_left_in[200]}),
		.sram(mux_2level_tapbuf_size18_9_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_9_sram_inv[0:9]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size18 mux_top_track_200 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[34], chanx_right_in[107], chanx_right_in[112], chanx_right_in[189], chanx_left_in[44], chanx_left_in[121], chanx_left_in[135], chanx_left_in[198]}),
		.sram(mux_2level_tapbuf_size18_10_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_10_sram_inv[0:9]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size18 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[36], chanx_right_in[111], chanx_right_in[113], chanx_right_in[190], chanx_left_in[42], chanx_left_in[120], chanx_left_in[131], chanx_left_in[197]}),
		.sram(mux_2level_tapbuf_size18_11_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_11_sram_inv[0:9]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size18 mux_top_track_224 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[38], chanx_right_in[116], chanx_right_in[119], chanx_right_in[193], chanx_left_in[40], chanx_left_in[117], chanx_left_in[123], chanx_left_in[194]}),
		.sram(mux_2level_tapbuf_size18_12_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_12_sram_inv[0:9]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size18 mux_top_track_232 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[40], chanx_right_in[117], chanx_right_in[123], chanx_right_in[194], chanx_left_in[38], chanx_left_in[116], chanx_left_in[119], chanx_left_in[193]}),
		.sram(mux_2level_tapbuf_size18_13_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_13_sram_inv[0:9]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size18 mux_top_track_240 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[41], chanx_right_in[118], chanx_right_in[127], chanx_right_in[196], chanx_left_in[37], chanx_left_in[114:115], chanx_left_in[192]}),
		.sram(mux_2level_tapbuf_size18_14_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_14_sram_inv[0:9]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size18 mux_top_track_248 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[42], chanx_right_in[120], chanx_right_in[131], chanx_right_in[197], chanx_left_in[36], chanx_left_in[111], chanx_left_in[113], chanx_left_in[190]}),
		.sram(mux_2level_tapbuf_size18_15_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_15_sram_inv[0:9]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size18 mux_top_track_256 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[44], chanx_right_in[121], chanx_right_in[135], chanx_right_in[198], chanx_left_in[34], chanx_left_in[107], chanx_left_in[112], chanx_left_in[189]}),
		.sram(mux_2level_tapbuf_size18_16_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_16_sram_inv[0:9]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size18 mux_top_track_264 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[45], chanx_right_in[122], chanx_right_in[139], chanx_right_in[200], chanx_left_in[33], chanx_left_in[103], chanx_left_in[110], chanx_left_in[188]}),
		.sram(mux_2level_tapbuf_size18_17_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_17_sram_inv[0:9]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size18 mux_top_track_272 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[46], chanx_right_in[124], chanx_right_in[143], chanx_right_in[201], chanx_left_in[32], chanx_left_in[99], chanx_left_in[109], chanx_left_in[186]}),
		.sram(mux_2level_tapbuf_size18_18_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_18_sram_inv[0:9]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size18 mux_top_track_280 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[48], chanx_right_in[125], chanx_right_in[147], chanx_right_in[202], chanx_left_in[30], chanx_left_in[95], chanx_left_in[108], chanx_left_in[185]}),
		.sram(mux_2level_tapbuf_size18_19_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_19_sram_inv[0:9]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size18 mux_top_track_296 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[50], chanx_right_in[128], chanx_right_in[155], chanx_right_in[205], chanx_left_in[28], chanx_left_in[87], chanx_left_in[105], chanx_left_in[182]}),
		.sram(mux_2level_tapbuf_size18_20_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_20_sram_inv[0:9]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size18 mux_top_track_304 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[52], chanx_right_in[129], chanx_right_in[159], chanx_right_in[206], chanx_left_in[26], chanx_left_in[83], chanx_left_in[104], chanx_left_in[181]}),
		.sram(mux_2level_tapbuf_size18_21_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_21_sram_inv[0:9]),
		.out(chany_top_out[152]));

	mux_2level_tapbuf_size18 mux_top_track_312 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[53], chanx_right_in[130], chanx_right_in[163], chanx_right_in[208], chanx_left_in[25], chanx_left_in[79], chanx_left_in[102], chanx_left_in[180]}),
		.sram(mux_2level_tapbuf_size18_22_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_22_sram_inv[0:9]),
		.out(chany_top_out[156]));

	mux_2level_tapbuf_size18 mux_top_track_320 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[54], chanx_right_in[132], chanx_right_in[167], chanx_right_in[209], chanx_left_in[24], chanx_left_in[75], chanx_left_in[101], chanx_left_in[178]}),
		.sram(mux_2level_tapbuf_size18_23_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_23_sram_inv[0:9]),
		.out(chany_top_out[160]));

	mux_2level_tapbuf_size18 mux_top_track_328 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[56], chanx_right_in[133], chanx_right_in[171], chanx_right_in[210], chanx_left_in[22], chanx_left_in[71], chanx_left_in[100], chanx_left_in[177]}),
		.sram(mux_2level_tapbuf_size18_24_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_24_sram_inv[0:9]),
		.out(chany_top_out[164]));

	mux_2level_tapbuf_size18 mux_top_track_336 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[57], chanx_right_in[134], chanx_right_in[175], chanx_right_in[212], chanx_left_in[21], chanx_left_in[67], chanx_left_in[98], chanx_left_in[176]}),
		.sram(mux_2level_tapbuf_size18_25_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_25_sram_inv[0:9]),
		.out(chany_top_out[168]));

	mux_2level_tapbuf_size18 mux_top_track_344 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[58], chanx_right_in[136], chanx_right_in[179], chanx_right_in[213], chanx_left_in[20], chanx_left_in[63], chanx_left_in[97], chanx_left_in[174]}),
		.sram(mux_2level_tapbuf_size18_26_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_26_sram_inv[0:9]),
		.out(chany_top_out[172]));

	mux_2level_tapbuf_size18 mux_top_track_352 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[60], chanx_right_in[137], chanx_right_in[183], chanx_right_in[214], chanx_left_in[18], chanx_left_in[59], chanx_left_in[96], chanx_left_in[173]}),
		.sram(mux_2level_tapbuf_size18_27_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_27_sram_inv[0:9]),
		.out(chany_top_out[176]));

	mux_2level_tapbuf_size18 mux_top_track_368 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[62], chanx_right_in[140], chanx_right_in[191], chanx_right_in[217], chanx_left_in[16], chanx_left_in[51], chanx_left_in[93], chanx_left_in[170]}),
		.sram(mux_2level_tapbuf_size18_28_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_28_sram_inv[0:9]),
		.out(chany_top_out[184]));

	mux_2level_tapbuf_size18 mux_top_track_376 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[64], chanx_right_in[141], chanx_right_in[195], chanx_right_in[218], chanx_left_in[14], chanx_left_in[47], chanx_left_in[92], chanx_left_in[169]}),
		.sram(mux_2level_tapbuf_size18_29_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_29_sram_inv[0:9]),
		.out(chany_top_out[188]));

	mux_2level_tapbuf_size18 mux_top_track_384 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[65], chanx_right_in[142], chanx_right_in[199], chanx_right_in[220], chanx_left_in[13], chanx_left_in[43], chanx_left_in[90], chanx_left_in[168]}),
		.sram(mux_2level_tapbuf_size18_30_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_30_sram_inv[0:9]),
		.out(chany_top_out[192]));

	mux_2level_tapbuf_size18 mux_top_track_392 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_, chanx_right_in[66], chanx_right_in[144], chanx_right_in[203], chanx_right_in[221], chanx_left_in[12], chanx_left_in[39], chanx_left_in[89], chanx_left_in[166]}),
		.sram(mux_2level_tapbuf_size18_31_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_31_sram_inv[0:9]),
		.out(chany_top_out[196]));

	mux_2level_tapbuf_size18 mux_top_track_400 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_, chanx_right_in[68], chanx_right_in[145], chanx_right_in[207], chanx_right_in[222], chanx_left_in[10], chanx_left_in[35], chanx_left_in[88], chanx_left_in[165]}),
		.sram(mux_2level_tapbuf_size18_32_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_32_sram_inv[0:9]),
		.out(chany_top_out[200]));

	mux_2level_tapbuf_size18 mux_top_track_408 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_, chanx_right_in[69], chanx_right_in[146], chanx_right_in[211], chanx_right_in[224], chanx_left_in[9], chanx_left_in[31], chanx_left_in[86], chanx_left_in[164]}),
		.sram(mux_2level_tapbuf_size18_33_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_33_sram_inv[0:9]),
		.out(chany_top_out[204]));

	mux_2level_tapbuf_size18 mux_top_track_416 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_, chanx_right_in[70], chanx_right_in[148], chanx_right_in[215], chanx_right_in[225], chanx_left_in[8], chanx_left_in[27], chanx_left_in[85], chanx_left_in[162]}),
		.sram(mux_2level_tapbuf_size18_34_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_34_sram_inv[0:9]),
		.out(chany_top_out[208]));

	mux_2level_tapbuf_size18 mux_top_track_424 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[72], chanx_right_in[149], chanx_right_in[219], chanx_right_in[226], chanx_left_in[6], chanx_left_in[23], chanx_left_in[84], chanx_left_in[161]}),
		.sram(mux_2level_tapbuf_size18_35_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_35_sram_inv[0:9]),
		.out(chany_top_out[212]));

	mux_2level_tapbuf_size18 mux_top_track_432 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_, chanx_right_in[73], chanx_right_in[150], chanx_right_in[223], chanx_left_in[5], chanx_left_in[19], chanx_left_in[82], chanx_left_in[160]}),
		.sram(mux_2level_tapbuf_size18_36_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_36_sram_inv[0:9]),
		.out(chany_top_out[216]));

	mux_2level_tapbuf_size18 mux_top_track_456 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_, chanx_right_in[0], chanx_right_in[3], chanx_right_in[77], chanx_right_in[154], chanx_left_in[1], chanx_left_in[7], chanx_left_in[78], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size18_37_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size18_37_sram_inv[0:9]),
		.out(chany_top_out[228]));

	mux_2level_tapbuf_size18_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_0_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_1_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_2_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_2_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_3_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_3_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_4_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_4_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_5_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_5_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_6_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_6_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_7_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_7_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_8_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_8_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_9_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_9_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_10_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_10_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_11_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_11_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_12_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_12_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_13_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_13_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_14_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_14_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_15_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_15_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_16_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_16_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_17_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_17_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_18_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_18_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_19_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_19_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_20_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_20_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_21_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_21_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_22_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_22_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_23_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_23_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_24_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_24_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_25_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_25_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_26_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_26_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_27_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_27_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size19_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_28_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_28_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_376 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_29_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_29_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_30_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_30_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_31_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_31_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_32_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_32_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_33_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_33_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_34_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_34_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_35_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_35_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_432 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_36_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_36_sram_inv[0:9]));

	mux_2level_tapbuf_size18_mem mem_top_track_456 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size17_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size18_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size18_37_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size18_37_sram_inv[0:9]));

	mux_2level_tapbuf_size17 mux_top_track_440 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_, chanx_right_in[74], chanx_right_in[152], chanx_right_in[227], chanx_left_in[4], chanx_left_in[15], chanx_left_in[81], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size17_0_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size17_0_sram_inv[0:9]),
		.out(chany_top_out[220]));

	mux_2level_tapbuf_size17 mux_top_track_448 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[76], chanx_right_in[153], chanx_right_in[228], chanx_left_in[2], chanx_left_in[11], chanx_left_in[80], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size17_1_sram[0:9]),
		.sram_inv(mux_2level_tapbuf_size17_1_sram_inv[0:9]),
		.out(chany_top_out[224]));

	mux_2level_tapbuf_size17_mem mem_top_track_440 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size17_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size17_0_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size17_0_sram_inv[0:9]));

	mux_2level_tapbuf_size17_mem mem_top_track_448 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size17_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size17_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size17_1_sram[0:9]),
		.mem_outb(mux_2level_tapbuf_size17_1_sram_inv[0:9]));

	mux_2level_tapbuf_size12 mux_right_track_0 (
		.in({chany_top_in[76], chany_top_in[153], chany_top_in[228], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[74], chany_bottom_in[152], chany_bottom_in[227]}),
		.sram(mux_2level_tapbuf_size12_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_0_sram_inv[0:7]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size12_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size18_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_0_sram_inv[0:7]));

	mux_2level_tapbuf_size13 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[77], chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[73], chany_bottom_in[150], chany_bottom_in[223]}),
		.sram(mux_2level_tapbuf_size13_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_0_sram_inv[0:7]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size13 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[86], chany_top_in[164], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[64], chany_bottom_in[141], chany_bottom_in[195], chany_bottom_in[218]}),
		.sram(mux_2level_tapbuf_size13_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_1_sram_inv[0:7]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size13 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[98], chany_top_in[176], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[52], chany_bottom_in[129], chany_bottom_in[159], chany_bottom_in[206]}),
		.sram(mux_2level_tapbuf_size13_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_2_sram_inv[0:7]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size13 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[103], chany_top_in[110], chany_top_in[188], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[40], chany_bottom_in[117], chany_bottom_in[123], chany_bottom_in[194]}),
		.sram(mux_2level_tapbuf_size13_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_3_sram_inv[0:7]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size13 mux_right_track_280 (
		.in({chany_top_in[45], chany_top_in[122], chany_top_in[139], chany_top_in[200], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[105], chany_bottom_in[182]}),
		.sram(mux_2level_tapbuf_size13_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_4_sram_inv[0:7]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size13 mux_right_track_352 (
		.in({chany_top_in[57], chany_top_in[134], chany_top_in[175], chany_top_in[212], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[93], chany_bottom_in[170]}),
		.sram(mux_2level_tapbuf_size13_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_5_sram_inv[0:7]),
		.out(chanx_right_out[176]));

	mux_2level_tapbuf_size13 mux_right_track_384 (
		.in({chany_top_in[62], chany_top_in[140], chany_top_in[191], chany_top_in[217], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[88], chany_bottom_in[165]}),
		.sram(mux_2level_tapbuf_size13_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_6_sram_inv[0:7]),
		.out(chanx_right_out[192]));

	mux_2level_tapbuf_size13 mux_right_track_392 (
		.in({chany_top_in[64], chany_top_in[141], chany_top_in[195], chany_top_in[218], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[86], chany_bottom_in[164]}),
		.sram(mux_2level_tapbuf_size13_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_7_sram_inv[0:7]),
		.out(chanx_right_out[196]));

	mux_2level_tapbuf_size13 mux_right_track_400 (
		.in({chany_top_in[65], chany_top_in[142], chany_top_in[199], chany_top_in[220], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[85], chany_bottom_in[162]}),
		.sram(mux_2level_tapbuf_size13_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_8_sram_inv[0:7]),
		.out(chanx_right_out[200]));

	mux_2level_tapbuf_size13 mux_right_track_408 (
		.in({chany_top_in[66], chany_top_in[144], chany_top_in[203], chany_top_in[221], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[84], chany_bottom_in[161]}),
		.sram(mux_2level_tapbuf_size13_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_9_sram_inv[0:7]),
		.out(chanx_right_out[204]));

	mux_2level_tapbuf_size13 mux_right_track_416 (
		.in({chany_top_in[68], chany_top_in[145], chany_top_in[207], chany_top_in[222], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[82], chany_bottom_in[160]}),
		.sram(mux_2level_tapbuf_size13_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_10_sram_inv[0:7]),
		.out(chanx_right_out[208]));

	mux_2level_tapbuf_size13 mux_right_track_424 (
		.in({chany_top_in[69], chany_top_in[146], chany_top_in[211], chany_top_in[224], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[81], chany_bottom_in[158]}),
		.sram(mux_2level_tapbuf_size13_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_11_sram_inv[0:7]),
		.out(chanx_right_out[212]));

	mux_2level_tapbuf_size13 mux_right_track_448 (
		.in({chany_top_in[73], chany_top_in[150], chany_top_in[223], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[77], chany_bottom_in[154]}),
		.sram(mux_2level_tapbuf_size13_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_12_sram_inv[0:7]),
		.out(chanx_right_out[224]));

	mux_2level_tapbuf_size13_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_0_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_1_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_2_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_3_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_4_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_5_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_6_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_7_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_8_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_9_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_10_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_11_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_448 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_12_sram_inv[0:7]));

	mux_2level_tapbuf_size14 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[78], chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[72], chany_bottom_in[149], chany_bottom_in[219], chany_bottom_in[226]}),
		.sram(mux_2level_tapbuf_size14_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_0_sram_inv[0:7]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size14 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[80], chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[70], chany_bottom_in[148], chany_bottom_in[215], chany_bottom_in[225]}),
		.sram(mux_2level_tapbuf_size14_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_1_sram_inv[0:7]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size14 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[81], chany_top_in[158], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[69], chany_bottom_in[146], chany_bottom_in[211], chany_bottom_in[224]}),
		.sram(mux_2level_tapbuf_size14_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_2_sram_inv[0:7]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size14 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[82], chany_top_in[160], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[68], chany_bottom_in[145], chany_bottom_in[207], chany_bottom_in[222]}),
		.sram(mux_2level_tapbuf_size14_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_3_sram_inv[0:7]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size14 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[84], chany_top_in[161], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[66], chany_bottom_in[144], chany_bottom_in[203], chany_bottom_in[221]}),
		.sram(mux_2level_tapbuf_size14_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_4_sram_inv[0:7]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size14 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[85], chany_top_in[162], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[65], chany_bottom_in[142], chany_bottom_in[199], chany_bottom_in[220]}),
		.sram(mux_2level_tapbuf_size14_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_5_sram_inv[0:7]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size14 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[88], chany_top_in[165], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[62], chany_bottom_in[140], chany_bottom_in[191], chany_bottom_in[217]}),
		.sram(mux_2level_tapbuf_size14_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_6_sram_inv[0:7]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size14 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[89], chany_top_in[166], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[61], chany_bottom_in[138], chany_bottom_in[187], chany_bottom_in[216]}),
		.sram(mux_2level_tapbuf_size14_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_7_sram_inv[0:7]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size14 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[90], chany_top_in[168], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[60], chany_bottom_in[137], chany_bottom_in[183], chany_bottom_in[214]}),
		.sram(mux_2level_tapbuf_size14_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_8_sram_inv[0:7]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size14 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[92], chany_top_in[169], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[58], chany_bottom_in[136], chany_bottom_in[179], chany_bottom_in[213]}),
		.sram(mux_2level_tapbuf_size14_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_9_sram_inv[0:7]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size14 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[93], chany_top_in[170], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[57], chany_bottom_in[134], chany_bottom_in[175], chany_bottom_in[212]}),
		.sram(mux_2level_tapbuf_size14_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_10_sram_inv[0:7]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size14 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[94], chany_top_in[172], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[56], chany_bottom_in[133], chany_bottom_in[171], chany_bottom_in[210]}),
		.sram(mux_2level_tapbuf_size14_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_11_sram_inv[0:7]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size14 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[96], chany_top_in[173], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[54], chany_bottom_in[132], chany_bottom_in[167], chany_bottom_in[209]}),
		.sram(mux_2level_tapbuf_size14_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_12_sram_inv[0:7]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size14 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[97], chany_top_in[174], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[53], chany_bottom_in[130], chany_bottom_in[163], chany_bottom_in[208]}),
		.sram(mux_2level_tapbuf_size14_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_13_sram_inv[0:7]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size14 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[100], chany_top_in[177], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[50], chany_bottom_in[128], chany_bottom_in[155], chany_bottom_in[205]}),
		.sram(mux_2level_tapbuf_size14_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_14_sram_inv[0:7]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size14 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[101], chany_top_in[178], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[49], chany_bottom_in[126], chany_bottom_in[151], chany_bottom_in[204]}),
		.sram(mux_2level_tapbuf_size14_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_15_sram_inv[0:7]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size14 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[102], chany_top_in[180], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[48], chany_bottom_in[125], chany_bottom_in[147], chany_bottom_in[202]}),
		.sram(mux_2level_tapbuf_size14_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_16_sram_inv[0:7]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size14 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[104], chany_top_in[181], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[46], chany_bottom_in[124], chany_bottom_in[143], chany_bottom_in[201]}),
		.sram(mux_2level_tapbuf_size14_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_17_sram_inv[0:7]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size14 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[105], chany_top_in[182], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[45], chany_bottom_in[122], chany_bottom_in[139], chany_bottom_in[200]}),
		.sram(mux_2level_tapbuf_size14_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_18_sram_inv[0:7]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size14 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[106], chany_top_in[184], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[44], chany_bottom_in[121], chany_bottom_in[135], chany_bottom_in[198]}),
		.sram(mux_2level_tapbuf_size14_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_19_sram_inv[0:7]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size14 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[95], chany_top_in[108], chany_top_in[185], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[42], chany_bottom_in[120], chany_bottom_in[131], chany_bottom_in[197]}),
		.sram(mux_2level_tapbuf_size14_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_20_sram_inv[0:7]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size14 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[99], chany_top_in[109], chany_top_in[186], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[41], chany_bottom_in[118], chany_bottom_in[127], chany_bottom_in[196]}),
		.sram(mux_2level_tapbuf_size14_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_21_sram_inv[0:7]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size14 mux_right_track_216 (
		.in({chany_top_in[34], chany_top_in[107], chany_top_in[112], chany_top_in[189], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[38], chany_bottom_in[116], chany_bottom_in[119], chany_bottom_in[193]}),
		.sram(mux_2level_tapbuf_size14_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_22_sram_inv[0:7]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size14 mux_right_track_224 (
		.in({chany_top_in[36], chany_top_in[111], chany_top_in[113], chany_top_in[190], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[37], chany_bottom_in[114:115], chany_bottom_in[192]}),
		.sram(mux_2level_tapbuf_size14_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_23_sram_inv[0:7]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size14 mux_right_track_232 (
		.in({chany_top_in[37], chany_top_in[114:115], chany_top_in[192], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[36], chany_bottom_in[111], chany_bottom_in[113], chany_bottom_in[190]}),
		.sram(mux_2level_tapbuf_size14_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_24_sram_inv[0:7]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size14 mux_right_track_240 (
		.in({chany_top_in[38], chany_top_in[116], chany_top_in[119], chany_top_in[193], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[34], chany_bottom_in[107], chany_bottom_in[112], chany_bottom_in[189]}),
		.sram(mux_2level_tapbuf_size14_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_25_sram_inv[0:7]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size14 mux_right_track_248 (
		.in({chany_top_in[40], chany_top_in[117], chany_top_in[123], chany_top_in[194], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[33], chany_bottom_in[103], chany_bottom_in[110], chany_bottom_in[188]}),
		.sram(mux_2level_tapbuf_size14_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_26_sram_inv[0:7]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size14 mux_right_track_256 (
		.in({chany_top_in[41], chany_top_in[118], chany_top_in[127], chany_top_in[196], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[32], chany_bottom_in[99], chany_bottom_in[109], chany_bottom_in[186]}),
		.sram(mux_2level_tapbuf_size14_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_27_sram_inv[0:7]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size14 mux_right_track_264 (
		.in({chany_top_in[42], chany_top_in[120], chany_top_in[131], chany_top_in[197], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[30], chany_bottom_in[95], chany_bottom_in[108], chany_bottom_in[185]}),
		.sram(mux_2level_tapbuf_size14_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_28_sram_inv[0:7]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size14 mux_right_track_272 (
		.in({chany_top_in[44], chany_top_in[121], chany_top_in[135], chany_top_in[198], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[106], chany_bottom_in[184]}),
		.sram(mux_2level_tapbuf_size14_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_29_sram_inv[0:7]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size14 mux_right_track_288 (
		.in({chany_top_in[46], chany_top_in[124], chany_top_in[143], chany_top_in[201], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[104], chany_bottom_in[181]}),
		.sram(mux_2level_tapbuf_size14_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_30_sram_inv[0:7]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size14 mux_right_track_296 (
		.in({chany_top_in[48], chany_top_in[125], chany_top_in[147], chany_top_in[202], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[102], chany_bottom_in[180]}),
		.sram(mux_2level_tapbuf_size14_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_31_sram_inv[0:7]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size14 mux_right_track_304 (
		.in({chany_top_in[49], chany_top_in[126], chany_top_in[151], chany_top_in[204], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[101], chany_bottom_in[178]}),
		.sram(mux_2level_tapbuf_size14_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_32_sram_inv[0:7]),
		.out(chanx_right_out[152]));

	mux_2level_tapbuf_size14 mux_right_track_312 (
		.in({chany_top_in[50], chany_top_in[128], chany_top_in[155], chany_top_in[205], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[100], chany_bottom_in[177]}),
		.sram(mux_2level_tapbuf_size14_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_33_sram_inv[0:7]),
		.out(chanx_right_out[156]));

	mux_2level_tapbuf_size14 mux_right_track_320 (
		.in({chany_top_in[52], chany_top_in[129], chany_top_in[159], chany_top_in[206], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[98], chany_bottom_in[176]}),
		.sram(mux_2level_tapbuf_size14_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_34_sram_inv[0:7]),
		.out(chanx_right_out[160]));

	mux_2level_tapbuf_size14 mux_right_track_328 (
		.in({chany_top_in[53], chany_top_in[130], chany_top_in[163], chany_top_in[208], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[97], chany_bottom_in[174]}),
		.sram(mux_2level_tapbuf_size14_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_35_sram_inv[0:7]),
		.out(chanx_right_out[164]));

	mux_2level_tapbuf_size14 mux_right_track_336 (
		.in({chany_top_in[54], chany_top_in[132], chany_top_in[167], chany_top_in[209], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[96], chany_bottom_in[173]}),
		.sram(mux_2level_tapbuf_size14_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_36_sram_inv[0:7]),
		.out(chanx_right_out[168]));

	mux_2level_tapbuf_size14 mux_right_track_344 (
		.in({chany_top_in[56], chany_top_in[133], chany_top_in[171], chany_top_in[210], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[94], chany_bottom_in[172]}),
		.sram(mux_2level_tapbuf_size14_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_37_sram_inv[0:7]),
		.out(chanx_right_out[172]));

	mux_2level_tapbuf_size14 mux_right_track_360 (
		.in({chany_top_in[58], chany_top_in[136], chany_top_in[179], chany_top_in[213], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[92], chany_bottom_in[169]}),
		.sram(mux_2level_tapbuf_size14_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_38_sram_inv[0:7]),
		.out(chanx_right_out[180]));

	mux_2level_tapbuf_size14 mux_right_track_368 (
		.in({chany_top_in[60], chany_top_in[137], chany_top_in[183], chany_top_in[214], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[90], chany_bottom_in[168]}),
		.sram(mux_2level_tapbuf_size14_39_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_39_sram_inv[0:7]),
		.out(chanx_right_out[184]));

	mux_2level_tapbuf_size14 mux_right_track_376 (
		.in({chany_top_in[61], chany_top_in[138], chany_top_in[187], chany_top_in[216], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[89], chany_bottom_in[166]}),
		.sram(mux_2level_tapbuf_size14_40_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_40_sram_inv[0:7]),
		.out(chanx_right_out[188]));

	mux_2level_tapbuf_size14 mux_right_track_432 (
		.in({chany_top_in[70], chany_top_in[148], chany_top_in[215], chany_top_in[225], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[80], chany_bottom_in[157]}),
		.sram(mux_2level_tapbuf_size14_41_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_41_sram_inv[0:7]),
		.out(chanx_right_out[216]));

	mux_2level_tapbuf_size14 mux_right_track_440 (
		.in({chany_top_in[72], chany_top_in[149], chany_top_in[219], chany_top_in[226], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[78], chany_bottom_in[156]}),
		.sram(mux_2level_tapbuf_size14_42_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_42_sram_inv[0:7]),
		.out(chanx_right_out[220]));

	mux_2level_tapbuf_size14_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_0_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_1_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_2_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_3_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_4_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_5_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_6_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_7_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_8_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_9_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_10_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_11_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_12_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_13_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_14_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_15_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_16_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_17_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_18_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_19_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_20_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_21_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_22_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_23_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_24_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_25_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_26_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_27_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_28_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_29_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_30_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_31_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_32_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_33_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_34_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_35_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_36_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_37_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_38_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_39_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_39_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_376 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_40_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_40_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_432 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_41_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_41_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_right_track_440 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_42_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_42_sram_inv[0:7]));

	mux_2level_tapbuf_size11 mux_right_track_456 (
		.in({chany_top_in[74], chany_top_in[152], chany_top_in[227], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, chany_bottom_in[76], chany_bottom_in[153], chany_bottom_in[228]}),
		.sram(mux_2level_tapbuf_size11_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_0_sram_inv[0:7]),
		.out(chanx_right_out[228]));

	mux_2level_tapbuf_size11_mem mem_right_track_456 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_0_sram_inv[0:7]));

	mux_2level_tapbuf_size9 mux_bottom_track_1 (
		.in({chanx_right_in[74], chanx_right_in[152], chanx_right_in[227], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[1], chanx_left_in[7], chanx_left_in[78], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size9_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_0_sram_inv[0:7]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size9 mux_bottom_track_9 (
		.in({chanx_right_in[73], chanx_right_in[150], chanx_right_in[223], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[2], chanx_left_in[11], chanx_left_in[80], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size9_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_1_sram_inv[0:7]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size9 mux_bottom_track_49 (
		.in({chanx_right_in[66], chanx_right_in[144], chanx_right_in[203], chanx_right_in[221], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[9], chanx_left_in[31], chanx_left_in[86], chanx_left_in[164]}),
		.sram(mux_2level_tapbuf_size9_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_2_sram_inv[0:7]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size9 mux_bottom_track_57 (
		.in({chanx_right_in[65], chanx_right_in[142], chanx_right_in[199], chanx_right_in[220], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[10], chanx_left_in[35], chanx_left_in[88], chanx_left_in[165]}),
		.sram(mux_2level_tapbuf_size9_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_3_sram_inv[0:7]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size9 mux_bottom_track_65 (
		.in({chanx_right_in[64], chanx_right_in[141], chanx_right_in[195], chanx_right_in[218], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[12], chanx_left_in[39], chanx_left_in[89], chanx_left_in[166]}),
		.sram(mux_2level_tapbuf_size9_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_4_sram_inv[0:7]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size9 mux_bottom_track_81 (
		.in({chanx_right_in[61], chanx_right_in[138], chanx_right_in[187], chanx_right_in[216], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[14], chanx_left_in[47], chanx_left_in[92], chanx_left_in[169]}),
		.sram(mux_2level_tapbuf_size9_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_5_sram_inv[0:7]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size9 mux_bottom_track_89 (
		.in({chanx_right_in[60], chanx_right_in[137], chanx_right_in[183], chanx_right_in[214], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[16], chanx_left_in[51], chanx_left_in[93], chanx_left_in[170]}),
		.sram(mux_2level_tapbuf_size9_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_6_sram_inv[0:7]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size9 mux_bottom_track_97 (
		.in({chanx_right_in[58], chanx_right_in[136], chanx_right_in[179], chanx_right_in[213], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[17], chanx_left_in[55], chanx_left_in[94], chanx_left_in[172]}),
		.sram(mux_2level_tapbuf_size9_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_7_sram_inv[0:7]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size9 mux_bottom_track_105 (
		.in({chanx_right_in[57], chanx_right_in[134], chanx_right_in[175], chanx_right_in[212], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[18], chanx_left_in[59], chanx_left_in[96], chanx_left_in[173]}),
		.sram(mux_2level_tapbuf_size9_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_8_sram_inv[0:7]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size9 mux_bottom_track_113 (
		.in({chanx_right_in[56], chanx_right_in[133], chanx_right_in[171], chanx_right_in[210], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[20], chanx_left_in[63], chanx_left_in[97], chanx_left_in[174]}),
		.sram(mux_2level_tapbuf_size9_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_9_sram_inv[0:7]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size9 mux_bottom_track_121 (
		.in({chanx_right_in[54], chanx_right_in[132], chanx_right_in[167], chanx_right_in[209], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[21], chanx_left_in[67], chanx_left_in[98], chanx_left_in[176]}),
		.sram(mux_2level_tapbuf_size9_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_10_sram_inv[0:7]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size9 mux_bottom_track_129 (
		.in({chanx_right_in[53], chanx_right_in[130], chanx_right_in[163], chanx_right_in[208], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[22], chanx_left_in[71], chanx_left_in[100], chanx_left_in[177]}),
		.sram(mux_2level_tapbuf_size9_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_11_sram_inv[0:7]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size9 mux_bottom_track_137 (
		.in({chanx_right_in[52], chanx_right_in[129], chanx_right_in[159], chanx_right_in[206], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[24], chanx_left_in[75], chanx_left_in[101], chanx_left_in[178]}),
		.sram(mux_2level_tapbuf_size9_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_12_sram_inv[0:7]),
		.out(chany_bottom_out[68]));

	mux_2level_tapbuf_size9 mux_bottom_track_153 (
		.in({chanx_right_in[49], chanx_right_in[126], chanx_right_in[151], chanx_right_in[204], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[26], chanx_left_in[83], chanx_left_in[104], chanx_left_in[181]}),
		.sram(mux_2level_tapbuf_size9_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_13_sram_inv[0:7]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size9 mux_bottom_track_161 (
		.in({chanx_right_in[48], chanx_right_in[125], chanx_right_in[147], chanx_right_in[202], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[28], chanx_left_in[87], chanx_left_in[105], chanx_left_in[182]}),
		.sram(mux_2level_tapbuf_size9_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_14_sram_inv[0:7]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size9 mux_bottom_track_169 (
		.in({chanx_right_in[46], chanx_right_in[124], chanx_right_in[143], chanx_right_in[201], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[29], chanx_left_in[91], chanx_left_in[106], chanx_left_in[184]}),
		.sram(mux_2level_tapbuf_size9_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_15_sram_inv[0:7]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size9 mux_bottom_track_177 (
		.in({chanx_right_in[45], chanx_right_in[122], chanx_right_in[139], chanx_right_in[200], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[30], chanx_left_in[95], chanx_left_in[108], chanx_left_in[185]}),
		.sram(mux_2level_tapbuf_size9_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_16_sram_inv[0:7]),
		.out(chany_bottom_out[88]));

	mux_2level_tapbuf_size9 mux_bottom_track_185 (
		.in({chanx_right_in[44], chanx_right_in[121], chanx_right_in[135], chanx_right_in[198], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[32], chanx_left_in[99], chanx_left_in[109], chanx_left_in[186]}),
		.sram(mux_2level_tapbuf_size9_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_17_sram_inv[0:7]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size9 mux_bottom_track_193 (
		.in({chanx_right_in[42], chanx_right_in[120], chanx_right_in[131], chanx_right_in[197], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[33], chanx_left_in[103], chanx_left_in[110], chanx_left_in[188]}),
		.sram(mux_2level_tapbuf_size9_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_18_sram_inv[0:7]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size9 mux_bottom_track_201 (
		.in({chanx_right_in[41], chanx_right_in[118], chanx_right_in[127], chanx_right_in[196], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[34], chanx_left_in[107], chanx_left_in[112], chanx_left_in[189]}),
		.sram(mux_2level_tapbuf_size9_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_19_sram_inv[0:7]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size9 mux_bottom_track_209 (
		.in({chanx_right_in[40], chanx_right_in[117], chanx_right_in[123], chanx_right_in[194], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[36], chanx_left_in[111], chanx_left_in[113], chanx_left_in[190]}),
		.sram(mux_2level_tapbuf_size9_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_20_sram_inv[0:7]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size9 mux_bottom_track_225 (
		.in({chanx_right_in[37], chanx_right_in[114:115], chanx_right_in[192], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[38], chanx_left_in[116], chanx_left_in[119], chanx_left_in[193]}),
		.sram(mux_2level_tapbuf_size9_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_21_sram_inv[0:7]),
		.out(chany_bottom_out[112]));

	mux_2level_tapbuf_size9 mux_bottom_track_233 (
		.in({chanx_right_in[36], chanx_right_in[111], chanx_right_in[113], chanx_right_in[190], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[40], chanx_left_in[117], chanx_left_in[123], chanx_left_in[194]}),
		.sram(mux_2level_tapbuf_size9_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_22_sram_inv[0:7]),
		.out(chany_bottom_out[116]));

	mux_2level_tapbuf_size9 mux_bottom_track_241 (
		.in({chanx_right_in[34], chanx_right_in[107], chanx_right_in[112], chanx_right_in[189], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[41], chanx_left_in[118], chanx_left_in[127], chanx_left_in[196]}),
		.sram(mux_2level_tapbuf_size9_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_23_sram_inv[0:7]),
		.out(chany_bottom_out[120]));

	mux_2level_tapbuf_size9 mux_bottom_track_249 (
		.in({chanx_right_in[33], chanx_right_in[103], chanx_right_in[110], chanx_right_in[188], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[42], chanx_left_in[120], chanx_left_in[131], chanx_left_in[197]}),
		.sram(mux_2level_tapbuf_size9_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_24_sram_inv[0:7]),
		.out(chany_bottom_out[124]));

	mux_2level_tapbuf_size9 mux_bottom_track_257 (
		.in({chanx_right_in[32], chanx_right_in[99], chanx_right_in[109], chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[44], chanx_left_in[121], chanx_left_in[135], chanx_left_in[198]}),
		.sram(mux_2level_tapbuf_size9_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_25_sram_inv[0:7]),
		.out(chany_bottom_out[128]));

	mux_2level_tapbuf_size9 mux_bottom_track_265 (
		.in({chanx_right_in[30], chanx_right_in[95], chanx_right_in[108], chanx_right_in[185], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[45], chanx_left_in[122], chanx_left_in[139], chanx_left_in[200]}),
		.sram(mux_2level_tapbuf_size9_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_26_sram_inv[0:7]),
		.out(chany_bottom_out[132]));

	mux_2level_tapbuf_size9 mux_bottom_track_273 (
		.in({chanx_right_in[29], chanx_right_in[91], chanx_right_in[106], chanx_right_in[184], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[46], chanx_left_in[124], chanx_left_in[143], chanx_left_in[201]}),
		.sram(mux_2level_tapbuf_size9_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_27_sram_inv[0:7]),
		.out(chany_bottom_out[136]));

	mux_2level_tapbuf_size9 mux_bottom_track_281 (
		.in({chanx_right_in[28], chanx_right_in[87], chanx_right_in[105], chanx_right_in[182], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[48], chanx_left_in[125], chanx_left_in[147], chanx_left_in[202]}),
		.sram(mux_2level_tapbuf_size9_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_28_sram_inv[0:7]),
		.out(chany_bottom_out[140]));

	mux_2level_tapbuf_size9 mux_bottom_track_297 (
		.in({chanx_right_in[25], chanx_right_in[79], chanx_right_in[102], chanx_right_in[180], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[50], chanx_left_in[128], chanx_left_in[155], chanx_left_in[205]}),
		.sram(mux_2level_tapbuf_size9_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_29_sram_inv[0:7]),
		.out(chany_bottom_out[148]));

	mux_2level_tapbuf_size9 mux_bottom_track_305 (
		.in({chanx_right_in[24], chanx_right_in[75], chanx_right_in[101], chanx_right_in[178], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[52], chanx_left_in[129], chanx_left_in[159], chanx_left_in[206]}),
		.sram(mux_2level_tapbuf_size9_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_30_sram_inv[0:7]),
		.out(chany_bottom_out[152]));

	mux_2level_tapbuf_size9 mux_bottom_track_313 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[100], chanx_right_in[177], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[53], chanx_left_in[130], chanx_left_in[163], chanx_left_in[208]}),
		.sram(mux_2level_tapbuf_size9_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_31_sram_inv[0:7]),
		.out(chany_bottom_out[156]));

	mux_2level_tapbuf_size9 mux_bottom_track_321 (
		.in({chanx_right_in[21], chanx_right_in[67], chanx_right_in[98], chanx_right_in[176], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[54], chanx_left_in[132], chanx_left_in[167], chanx_left_in[209]}),
		.sram(mux_2level_tapbuf_size9_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_32_sram_inv[0:7]),
		.out(chany_bottom_out[160]));

	mux_2level_tapbuf_size9 mux_bottom_track_329 (
		.in({chanx_right_in[20], chanx_right_in[63], chanx_right_in[97], chanx_right_in[174], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[56], chanx_left_in[133], chanx_left_in[171], chanx_left_in[210]}),
		.sram(mux_2level_tapbuf_size9_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_33_sram_inv[0:7]),
		.out(chany_bottom_out[164]));

	mux_2level_tapbuf_size9 mux_bottom_track_337 (
		.in({chanx_right_in[18], chanx_right_in[59], chanx_right_in[96], chanx_right_in[173], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[57], chanx_left_in[134], chanx_left_in[175], chanx_left_in[212]}),
		.sram(mux_2level_tapbuf_size9_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_34_sram_inv[0:7]),
		.out(chany_bottom_out[168]));

	mux_2level_tapbuf_size9 mux_bottom_track_345 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[94], chanx_right_in[172], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[58], chanx_left_in[136], chanx_left_in[179], chanx_left_in[213]}),
		.sram(mux_2level_tapbuf_size9_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_35_sram_inv[0:7]),
		.out(chany_bottom_out[172]));

	mux_2level_tapbuf_size9 mux_bottom_track_353 (
		.in({chanx_right_in[16], chanx_right_in[51], chanx_right_in[93], chanx_right_in[170], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[60], chanx_left_in[137], chanx_left_in[183], chanx_left_in[214]}),
		.sram(mux_2level_tapbuf_size9_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_36_sram_inv[0:7]),
		.out(chany_bottom_out[176]));

	mux_2level_tapbuf_size9 mux_bottom_track_369 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[90], chanx_right_in[168], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[62], chanx_left_in[140], chanx_left_in[191], chanx_left_in[217]}),
		.sram(mux_2level_tapbuf_size9_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_37_sram_inv[0:7]),
		.out(chany_bottom_out[184]));

	mux_2level_tapbuf_size9 mux_bottom_track_377 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[89], chanx_right_in[166], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[64], chanx_left_in[141], chanx_left_in[195], chanx_left_in[218]}),
		.sram(mux_2level_tapbuf_size9_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_38_sram_inv[0:7]),
		.out(chany_bottom_out[188]));

	mux_2level_tapbuf_size9 mux_bottom_track_385 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[88], chanx_right_in[165], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[65], chanx_left_in[142], chanx_left_in[199], chanx_left_in[220]}),
		.sram(mux_2level_tapbuf_size9_39_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_39_sram_inv[0:7]),
		.out(chany_bottom_out[192]));

	mux_2level_tapbuf_size9 mux_bottom_track_393 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[86], chanx_right_in[164], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[66], chanx_left_in[144], chanx_left_in[203], chanx_left_in[221]}),
		.sram(mux_2level_tapbuf_size9_40_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_40_sram_inv[0:7]),
		.out(chany_bottom_out[196]));

	mux_2level_tapbuf_size9 mux_bottom_track_401 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[85], chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[68], chanx_left_in[145], chanx_left_in[207], chanx_left_in[222]}),
		.sram(mux_2level_tapbuf_size9_41_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_41_sram_inv[0:7]),
		.out(chany_bottom_out[200]));

	mux_2level_tapbuf_size9 mux_bottom_track_409 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[84], chanx_right_in[161], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[69], chanx_left_in[146], chanx_left_in[211], chanx_left_in[224]}),
		.sram(mux_2level_tapbuf_size9_42_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_42_sram_inv[0:7]),
		.out(chany_bottom_out[204]));

	mux_2level_tapbuf_size9 mux_bottom_track_417 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[82], chanx_right_in[160], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[70], chanx_left_in[148], chanx_left_in[215], chanx_left_in[225]}),
		.sram(mux_2level_tapbuf_size9_43_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_43_sram_inv[0:7]),
		.out(chany_bottom_out[208]));

	mux_2level_tapbuf_size9 mux_bottom_track_425 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[81], chanx_right_in[158], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[72], chanx_left_in[149], chanx_left_in[219], chanx_left_in[226]}),
		.sram(mux_2level_tapbuf_size9_44_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_44_sram_inv[0:7]),
		.out(chany_bottom_out[212]));

	mux_2level_tapbuf_size9 mux_bottom_track_433 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[80], chanx_right_in[157], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[73], chanx_left_in[150], chanx_left_in[223]}),
		.sram(mux_2level_tapbuf_size9_45_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_45_sram_inv[0:7]),
		.out(chany_bottom_out[216]));

	mux_2level_tapbuf_size9 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[77], chany_top_in[154], chany_bottom_in[76], chany_bottom_in[153], chany_bottom_in[228], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_46_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_46_sram_inv[0:7]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size9 mux_left_track_33 (
		.in({chany_top_in[72], chany_top_in[149], chany_top_in[219], chany_top_in[226], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[81], chany_bottom_in[158], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_47_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_47_sram_inv[0:7]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size9 mux_left_track_73 (
		.in({chany_top_in[65], chany_top_in[142], chany_top_in[199], chany_top_in[220], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[88], chany_bottom_in[165], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_48_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_48_sram_inv[0:7]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size9 mux_left_track_81 (
		.in({chany_top_in[64], chany_top_in[141], chany_top_in[195], chany_top_in[218], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[89], chany_bottom_in[166], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_49_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_49_sram_inv[0:7]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size9 mux_left_track_89 (
		.in({chany_top_in[62], chany_top_in[140], chany_top_in[191], chany_top_in[217], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[90], chany_bottom_in[168], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size9_50_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_50_sram_inv[0:7]),
		.out(chanx_left_out[44]));

	mux_2level_tapbuf_size9 mux_left_track_97 (
		.in({chany_top_in[61], chany_top_in[138], chany_top_in[187], chany_top_in[216], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[92], chany_bottom_in[169], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size9_51_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_51_sram_inv[0:7]),
		.out(chanx_left_out[48]));

	mux_2level_tapbuf_size9 mux_left_track_105 (
		.in({chany_top_in[60], chany_top_in[137], chany_top_in[183], chany_top_in[214], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[93], chany_bottom_in[170], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_52_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_52_sram_inv[0:7]),
		.out(chanx_left_out[52]));

	mux_2level_tapbuf_size9 mux_left_track_145 (
		.in({chany_top_in[53], chany_top_in[130], chany_top_in[163], chany_top_in[208], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[100], chany_bottom_in[177], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_53_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_53_sram_inv[0:7]),
		.out(chanx_left_out[72]));

	mux_2level_tapbuf_size9 mux_left_track_153 (
		.in({chany_top_in[52], chany_top_in[129], chany_top_in[159], chany_top_in[206], chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[101], chany_bottom_in[178], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_54_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_54_sram_inv[0:7]),
		.out(chanx_left_out[76]));

	mux_2level_tapbuf_size9 mux_left_track_161 (
		.in({chany_top_in[50], chany_top_in[128], chany_top_in[155], chany_top_in[205], chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[102], chany_bottom_in[180], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size9_55_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_55_sram_inv[0:7]),
		.out(chanx_left_out[80]));

	mux_2level_tapbuf_size9 mux_left_track_169 (
		.in({chany_top_in[49], chany_top_in[126], chany_top_in[151], chany_top_in[204], chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[104], chany_bottom_in[181], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size9_56_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_56_sram_inv[0:7]),
		.out(chanx_left_out[84]));

	mux_2level_tapbuf_size9 mux_left_track_177 (
		.in({chany_top_in[48], chany_top_in[125], chany_top_in[147], chany_top_in[202], chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[105], chany_bottom_in[182], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_57_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_57_sram_inv[0:7]),
		.out(chanx_left_out[88]));

	mux_2level_tapbuf_size9 mux_left_track_217 (
		.in({chany_top_in[41], chany_top_in[118], chany_top_in[127], chany_top_in[196], chany_bottom_in[34], chany_bottom_in[107], chany_bottom_in[112], chany_bottom_in[189], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_58_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_58_sram_inv[0:7]),
		.out(chanx_left_out[108]));

	mux_2level_tapbuf_size9 mux_left_track_225 (
		.in({chany_top_in[40], chany_top_in[117], chany_top_in[123], chany_top_in[194], chany_bottom_in[36], chany_bottom_in[111], chany_bottom_in[113], chany_bottom_in[190], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_59_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_59_sram_inv[0:7]),
		.out(chanx_left_out[112]));

	mux_2level_tapbuf_size9 mux_left_track_233 (
		.in({chany_top_in[38], chany_top_in[116], chany_top_in[119], chany_top_in[193], chany_bottom_in[37], chany_bottom_in[114:115], chany_bottom_in[192], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size9_60_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_60_sram_inv[0:7]),
		.out(chanx_left_out[116]));

	mux_2level_tapbuf_size9 mux_left_track_241 (
		.in({chany_top_in[37], chany_top_in[114:115], chany_top_in[192], chany_bottom_in[38], chany_bottom_in[116], chany_bottom_in[119], chany_bottom_in[193], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size9_61_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_61_sram_inv[0:7]),
		.out(chanx_left_out[120]));

	mux_2level_tapbuf_size9 mux_left_track_249 (
		.in({chany_top_in[36], chany_top_in[111], chany_top_in[113], chany_top_in[190], chany_bottom_in[40], chany_bottom_in[117], chany_bottom_in[123], chany_bottom_in[194], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_62_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_62_sram_inv[0:7]),
		.out(chanx_left_out[124]));

	mux_2level_tapbuf_size9 mux_left_track_289 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[106], chany_top_in[184], chany_bottom_in[46], chany_bottom_in[124], chany_bottom_in[143], chany_bottom_in[201], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_63_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_63_sram_inv[0:7]),
		.out(chanx_left_out[144]));

	mux_2level_tapbuf_size9 mux_left_track_297 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[105], chany_top_in[182], chany_bottom_in[48], chany_bottom_in[125], chany_bottom_in[147], chany_bottom_in[202], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_64_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_64_sram_inv[0:7]),
		.out(chanx_left_out[148]));

	mux_2level_tapbuf_size9 mux_left_track_305 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[104], chany_top_in[181], chany_bottom_in[49], chany_bottom_in[126], chany_bottom_in[151], chany_bottom_in[204], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size9_65_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_65_sram_inv[0:7]),
		.out(chanx_left_out[152]));

	mux_2level_tapbuf_size9 mux_left_track_313 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[102], chany_top_in[180], chany_bottom_in[50], chany_bottom_in[128], chany_bottom_in[155], chany_bottom_in[205], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size9_66_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_66_sram_inv[0:7]),
		.out(chanx_left_out[156]));

	mux_2level_tapbuf_size9 mux_left_track_321 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[101], chany_top_in[178], chany_bottom_in[52], chany_bottom_in[129], chany_bottom_in[159], chany_bottom_in[206], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_67_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_67_sram_inv[0:7]),
		.out(chanx_left_out[160]));

	mux_2level_tapbuf_size9 mux_left_track_361 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[94], chany_top_in[172], chany_bottom_in[58], chany_bottom_in[136], chany_bottom_in[179], chany_bottom_in[213], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_68_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_68_sram_inv[0:7]),
		.out(chanx_left_out[180]));

	mux_2level_tapbuf_size9 mux_left_track_369 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[93], chany_top_in[170], chany_bottom_in[60], chany_bottom_in[137], chany_bottom_in[183], chany_bottom_in[214], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_69_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_69_sram_inv[0:7]),
		.out(chanx_left_out[184]));

	mux_2level_tapbuf_size9 mux_left_track_377 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[92], chany_top_in[169], chany_bottom_in[61], chany_bottom_in[138], chany_bottom_in[187], chany_bottom_in[216], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size9_70_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_70_sram_inv[0:7]),
		.out(chanx_left_out[188]));

	mux_2level_tapbuf_size9 mux_left_track_385 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[90], chany_top_in[168], chany_bottom_in[62], chany_bottom_in[140], chany_bottom_in[191], chany_bottom_in[217], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size9_71_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_71_sram_inv[0:7]),
		.out(chanx_left_out[192]));

	mux_2level_tapbuf_size9 mux_left_track_393 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[89], chany_top_in[166], chany_bottom_in[64], chany_bottom_in[141], chany_bottom_in[195], chany_bottom_in[218], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(mux_2level_tapbuf_size9_72_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_72_sram_inv[0:7]),
		.out(chanx_left_out[196]));

	mux_2level_tapbuf_size9 mux_left_track_433 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[82], chany_top_in[160], chany_bottom_in[70], chany_bottom_in[148], chany_bottom_in[215], chany_bottom_in[225], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_2level_tapbuf_size9_73_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_73_sram_inv[0:7]),
		.out(chanx_left_out[216]));

	mux_2level_tapbuf_size9 mux_left_track_441 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[81], chany_top_in[158], chany_bottom_in[72], chany_bottom_in[149], chany_bottom_in[219], chany_bottom_in[226], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size9_74_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_74_sram_inv[0:7]),
		.out(chanx_left_out[220]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_0_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_1_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_2_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_3_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_4_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_5_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_6_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_7_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_8_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_9_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_10_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_11_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_12_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_13_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_14_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_15_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_16_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_17_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_18_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_19_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_20_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_21_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_22_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_23_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_24_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_25_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_26_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_27_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_28_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_29_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_305 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_30_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_313 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_31_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_321 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_32_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_329 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_33_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_337 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_34_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_345 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_35_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_353 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_36_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_369 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_37_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_377 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_38_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_385 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_39_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_39_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_393 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_40_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_40_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_401 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_41_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_41_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_409 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_42_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_42_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_417 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_43_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_43_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_425 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_44_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_44_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_433 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_45_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_45_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_46_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_46_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_47_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_47_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_48_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_48_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_49_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_49_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_50_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_50_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_51_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_51_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_52_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_52_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_53_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_53_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_54_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_54_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_55_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_55_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_56_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_56_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_57_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_57_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_58_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_58_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_59_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_59_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_60_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_60_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_61_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_61_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_62_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_62_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_63_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_63_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_64_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_64_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_305 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_65_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_65_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_313 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_66_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_66_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_321 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_67_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_67_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_361 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_68_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_68_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_369 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_69_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_69_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_377 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_70_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_70_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_385 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_71_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_71_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_393 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_72_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_72_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_433 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_73_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_73_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_left_track_441 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_74_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_74_sram_inv[0:7]));

	mux_2level_tapbuf_size10 mux_bottom_track_17 (
		.in({chanx_right_in[72], chanx_right_in[149], chanx_right_in[219], chanx_right_in[226], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, chanx_left_in[4], chanx_left_in[15], chanx_left_in[81], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size10_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_0_sram_inv[0:7]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size10 mux_bottom_track_25 (
		.in({chanx_right_in[70], chanx_right_in[148], chanx_right_in[215], chanx_right_in[225], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[5], chanx_left_in[19], chanx_left_in[82], chanx_left_in[160]}),
		.sram(mux_2level_tapbuf_size10_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_1_sram_inv[0:7]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size10 mux_bottom_track_33 (
		.in({chanx_right_in[69], chanx_right_in[146], chanx_right_in[211], chanx_right_in[224], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[6], chanx_left_in[23], chanx_left_in[84], chanx_left_in[161]}),
		.sram(mux_2level_tapbuf_size10_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_2_sram_inv[0:7]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size10 mux_bottom_track_41 (
		.in({chanx_right_in[68], chanx_right_in[145], chanx_right_in[207], chanx_right_in[222], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[8], chanx_left_in[27], chanx_left_in[85], chanx_left_in[162]}),
		.sram(mux_2level_tapbuf_size10_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_3_sram_inv[0:7]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size10 mux_bottom_track_73 (
		.in({chanx_right_in[62], chanx_right_in[140], chanx_right_in[191], chanx_right_in[217], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[13], chanx_left_in[43], chanx_left_in[90], chanx_left_in[168]}),
		.sram(mux_2level_tapbuf_size10_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_4_sram_inv[0:7]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size10 mux_bottom_track_145 (
		.in({chanx_right_in[50], chanx_right_in[128], chanx_right_in[155], chanx_right_in[205], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[25], chanx_left_in[79], chanx_left_in[102], chanx_left_in[180]}),
		.sram(mux_2level_tapbuf_size10_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_5_sram_inv[0:7]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size10 mux_bottom_track_217 (
		.in({chanx_right_in[38], chanx_right_in[116], chanx_right_in[119], chanx_right_in[193], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[37], chanx_left_in[114:115], chanx_left_in[192]}),
		.sram(mux_2level_tapbuf_size10_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_6_sram_inv[0:7]),
		.out(chany_bottom_out[108]));

	mux_2level_tapbuf_size10 mux_bottom_track_289 (
		.in({chanx_right_in[26], chanx_right_in[83], chanx_right_in[104], chanx_right_in[181], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[49], chanx_left_in[126], chanx_left_in[151], chanx_left_in[204]}),
		.sram(mux_2level_tapbuf_size10_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_7_sram_inv[0:7]),
		.out(chany_bottom_out[144]));

	mux_2level_tapbuf_size10 mux_bottom_track_361 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[92], chanx_right_in[169], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[61], chanx_left_in[138], chanx_left_in[187], chanx_left_in[216]}),
		.sram(mux_2level_tapbuf_size10_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_8_sram_inv[0:7]),
		.out(chany_bottom_out[180]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_0_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_1_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_2_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_3_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_4_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_5_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_6_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_7_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_bottom_track_361 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_8_sram_inv[0:7]));

	mux_2level_tapbuf_size8 mux_bottom_track_441 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[78], chanx_right_in[156], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[74], chanx_left_in[152], chanx_left_in[227]}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chany_bottom_out[220]));

	mux_2level_tapbuf_size8 mux_bottom_track_449 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[77], chanx_right_in[154], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[76], chanx_left_in[153], chanx_left_in[228]}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chany_bottom_out[224]));

	mux_2level_tapbuf_size8 mux_bottom_track_457 (
		.in({chanx_right_in[76], chanx_right_in[153], chanx_right_in[228], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[0], chanx_left_in[3], chanx_left_in[77], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chany_bottom_out[228]));

	mux_2level_tapbuf_size8 mux_left_track_9 (
		.in({chany_top_in[76], chany_top_in[153], chany_top_in[228], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[77], chany_bottom_in[154], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size8 mux_left_track_17 (
		.in({chany_top_in[74], chany_top_in[152], chany_top_in[227], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[78], chany_bottom_in[156], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size8 mux_left_track_25 (
		.in({chany_top_in[73], chany_top_in[150], chany_top_in[223], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[80], chany_bottom_in[157], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size8 mux_left_track_41 (
		.in({chany_top_in[70], chany_top_in[148], chany_top_in[215], chany_top_in[225], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[82], chany_bottom_in[160]}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size8 mux_left_track_49 (
		.in({chany_top_in[69], chany_top_in[146], chany_top_in[211], chany_top_in[224], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[84], chany_bottom_in[161]}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size8 mux_left_track_57 (
		.in({chany_top_in[68], chany_top_in[145], chany_top_in[207], chany_top_in[222], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[85], chany_bottom_in[162]}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size8 mux_left_track_65 (
		.in({chany_top_in[66], chany_top_in[144], chany_top_in[203], chany_top_in[221], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[86], chany_bottom_in[164]}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size8 mux_left_track_113 (
		.in({chany_top_in[58], chany_top_in[136], chany_top_in[179], chany_top_in[213], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[94], chany_bottom_in[172]}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chanx_left_out[56]));

	mux_2level_tapbuf_size8 mux_left_track_121 (
		.in({chany_top_in[57], chany_top_in[134], chany_top_in[175], chany_top_in[212], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[96], chany_bottom_in[173]}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chanx_left_out[60]));

	mux_2level_tapbuf_size8 mux_left_track_129 (
		.in({chany_top_in[56], chany_top_in[133], chany_top_in[171], chany_top_in[210], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[97], chany_bottom_in[174]}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chanx_left_out[64]));

	mux_2level_tapbuf_size8 mux_left_track_137 (
		.in({chany_top_in[54], chany_top_in[132], chany_top_in[167], chany_top_in[209], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[98], chany_bottom_in[176]}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chanx_left_out[68]));

	mux_2level_tapbuf_size8 mux_left_track_185 (
		.in({chany_top_in[46], chany_top_in[124], chany_top_in[143], chany_top_in[201], chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[106], chany_bottom_in[184]}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chanx_left_out[92]));

	mux_2level_tapbuf_size8 mux_left_track_193 (
		.in({chany_top_in[45], chany_top_in[122], chany_top_in[139], chany_top_in[200], chany_bottom_in[30], chany_bottom_in[95], chany_bottom_in[108], chany_bottom_in[185]}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chanx_left_out[96]));

	mux_2level_tapbuf_size8 mux_left_track_201 (
		.in({chany_top_in[44], chany_top_in[121], chany_top_in[135], chany_top_in[198], chany_bottom_in[32], chany_bottom_in[99], chany_bottom_in[109], chany_bottom_in[186]}),
		.sram(mux_2level_tapbuf_size8_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_16_sram_inv[0:5]),
		.out(chanx_left_out[100]));

	mux_2level_tapbuf_size8 mux_left_track_209 (
		.in({chany_top_in[42], chany_top_in[120], chany_top_in[131], chany_top_in[197], chany_bottom_in[33], chany_bottom_in[103], chany_bottom_in[110], chany_bottom_in[188]}),
		.sram(mux_2level_tapbuf_size8_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_17_sram_inv[0:5]),
		.out(chanx_left_out[104]));

	mux_2level_tapbuf_size8 mux_left_track_257 (
		.in({chany_top_in[34], chany_top_in[107], chany_top_in[112], chany_top_in[189], chany_bottom_in[41], chany_bottom_in[118], chany_bottom_in[127], chany_bottom_in[196]}),
		.sram(mux_2level_tapbuf_size8_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_18_sram_inv[0:5]),
		.out(chanx_left_out[128]));

	mux_2level_tapbuf_size8 mux_left_track_265 (
		.in({chany_top_in[33], chany_top_in[103], chany_top_in[110], chany_top_in[188], chany_bottom_in[42], chany_bottom_in[120], chany_bottom_in[131], chany_bottom_in[197]}),
		.sram(mux_2level_tapbuf_size8_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_19_sram_inv[0:5]),
		.out(chanx_left_out[132]));

	mux_2level_tapbuf_size8 mux_left_track_273 (
		.in({chany_top_in[32], chany_top_in[99], chany_top_in[109], chany_top_in[186], chany_bottom_in[44], chany_bottom_in[121], chany_bottom_in[135], chany_bottom_in[198]}),
		.sram(mux_2level_tapbuf_size8_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_20_sram_inv[0:5]),
		.out(chanx_left_out[136]));

	mux_2level_tapbuf_size8 mux_left_track_281 (
		.in({chany_top_in[30], chany_top_in[95], chany_top_in[108], chany_top_in[185], chany_bottom_in[45], chany_bottom_in[122], chany_bottom_in[139], chany_bottom_in[200]}),
		.sram(mux_2level_tapbuf_size8_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_21_sram_inv[0:5]),
		.out(chanx_left_out[140]));

	mux_2level_tapbuf_size8 mux_left_track_329 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[100], chany_top_in[177], chany_bottom_in[53], chany_bottom_in[130], chany_bottom_in[163], chany_bottom_in[208]}),
		.sram(mux_2level_tapbuf_size8_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_22_sram_inv[0:5]),
		.out(chanx_left_out[164]));

	mux_2level_tapbuf_size8 mux_left_track_337 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[98], chany_top_in[176], chany_bottom_in[54], chany_bottom_in[132], chany_bottom_in[167], chany_bottom_in[209]}),
		.sram(mux_2level_tapbuf_size8_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_23_sram_inv[0:5]),
		.out(chanx_left_out[168]));

	mux_2level_tapbuf_size8 mux_left_track_345 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[97], chany_top_in[174], chany_bottom_in[56], chany_bottom_in[133], chany_bottom_in[171], chany_bottom_in[210]}),
		.sram(mux_2level_tapbuf_size8_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_24_sram_inv[0:5]),
		.out(chanx_left_out[172]));

	mux_2level_tapbuf_size8 mux_left_track_353 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[96], chany_top_in[173], chany_bottom_in[57], chany_bottom_in[134], chany_bottom_in[175], chany_bottom_in[212]}),
		.sram(mux_2level_tapbuf_size8_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_25_sram_inv[0:5]),
		.out(chanx_left_out[176]));

	mux_2level_tapbuf_size8 mux_left_track_401 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[88], chany_top_in[165], chany_bottom_in[65], chany_bottom_in[142], chany_bottom_in[199], chany_bottom_in[220]}),
		.sram(mux_2level_tapbuf_size8_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_26_sram_inv[0:5]),
		.out(chanx_left_out[200]));

	mux_2level_tapbuf_size8 mux_left_track_409 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[86], chany_top_in[164], chany_bottom_in[66], chany_bottom_in[144], chany_bottom_in[203], chany_bottom_in[221]}),
		.sram(mux_2level_tapbuf_size8_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_27_sram_inv[0:5]),
		.out(chanx_left_out[204]));

	mux_2level_tapbuf_size8 mux_left_track_417 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[85], chany_top_in[162], chany_bottom_in[68], chany_bottom_in[145], chany_bottom_in[207], chany_bottom_in[222]}),
		.sram(mux_2level_tapbuf_size8_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_28_sram_inv[0:5]),
		.out(chanx_left_out[208]));

	mux_2level_tapbuf_size8 mux_left_track_425 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[84], chany_top_in[161], chany_bottom_in[69], chany_bottom_in[146], chany_bottom_in[211], chany_bottom_in[224]}),
		.sram(mux_2level_tapbuf_size8_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_29_sram_inv[0:5]),
		.out(chanx_left_out[212]));

	mux_2level_tapbuf_size8 mux_left_track_449 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[80], chany_top_in[157], chany_bottom_in[73], chany_bottom_in[150], chany_bottom_in[223], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_2level_tapbuf_size8_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_30_sram_inv[0:5]),
		.out(chanx_left_out[224]));

	mux_2level_tapbuf_size8 mux_left_track_457 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[78], chany_top_in[156], chany_bottom_in[74], chany_bottom_in[152], chany_bottom_in[227], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(mux_2level_tapbuf_size8_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_31_sram_inv[0:5]),
		.out(chanx_left_out[228]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_441 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_449 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_457 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_16_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_17_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_18_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_19_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_20_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_21_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_329 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_22_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_337 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_23_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_345 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_24_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_353 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_25_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_401 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_26_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_409 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_27_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_417 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_28_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_425 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_29_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_449 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_30_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_left_track_457 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_31_sram_inv[0:5]));

endmodule
// ----- END Verilog module for sb_2__5_ -----

//----- Default net type -----
`default_nettype wire



