// localparams.sv
`ifndef localparamS_SV
`define localparamS_SV



// // Directories
// localparam string ROUTING_TABLES_DIR = 
//     (ROWS == 2 && COLUMNS == 2) ? "../routing_tables/mesh_2x2/" :
//     (ROWS == 3 && COLUMNS == 3) ? "../routing_tables/mesh_3x3/" :
//     (ROWS == 4 && COLUMNS == 4) ? "../routing_tables/mesh_4x4/" :
//     "../routing_tables/default/"; // Default this should be an error

`endif // localparamS_SV
