//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Formal Top-level netlist of Design: noc
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug  6 13:30:11 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module noc_top_formal_verification_random_tb;
// ----- Default clock port is added here since benchmark does not contain one -------
	reg [0:0] clk;

// ----- Shared inputs -------
	reg [0:0] n0_idata_p0_0_;
	reg [0:0] n0_idata_p0_1_;
	reg [0:0] n0_idata_p0_2_;
	reg [0:0] n0_idata_p0_3_;
	reg [0:0] n0_idata_p0_4_;
	reg [0:0] n0_idata_p0_5_;
	reg [0:0] n0_idata_p0_6_;
	reg [0:0] n0_idata_p0_7_;
	reg [0:0] n0_idata_p0_8_;
	reg [0:0] n0_idata_p0_9_;
	reg [0:0] n0_idata_p0_10_;
	reg [0:0] n0_idata_p0_11_;
	reg [0:0] n0_idata_p0_12_;
	reg [0:0] n0_idata_p0_13_;
	reg [0:0] n0_idata_p0_14_;
	reg [0:0] n0_idata_p0_15_;
	reg [0:0] n0_idata_p0_16_;
	reg [0:0] n0_idata_p0_17_;
	reg [0:0] n0_idata_p0_18_;
	reg [0:0] n0_idata_p0_19_;
	reg [0:0] n0_idata_p0_20_;
	reg [0:0] n0_idata_p0_21_;
	reg [0:0] n0_idata_p0_22_;
	reg [0:0] n0_idata_p0_23_;
	reg [0:0] n0_idata_p0_24_;
	reg [0:0] n0_idata_p0_25_;
	reg [0:0] n0_idata_p0_26_;
	reg [0:0] n0_idata_p0_27_;
	reg [0:0] n0_idata_p0_28_;
	reg [0:0] n0_idata_p0_29_;
	reg [0:0] n0_idata_p0_30_;
	reg [0:0] n0_idata_p0_31_;
	reg [0:0] n0_idata_p0_32_;
	reg [0:0] n0_idata_p0_33_;
	reg [0:0] n0_idata_p0_34_;
	reg [0:0] n0_ivalid_p0;
	reg [0:0] n0_ivch_p0;
	reg [0:0] n1_idata_p0_0_;
	reg [0:0] n1_idata_p0_1_;
	reg [0:0] n1_idata_p0_2_;
	reg [0:0] n1_idata_p0_3_;
	reg [0:0] n1_idata_p0_4_;
	reg [0:0] n1_idata_p0_5_;
	reg [0:0] n1_idata_p0_6_;
	reg [0:0] n1_idata_p0_7_;
	reg [0:0] n1_idata_p0_8_;
	reg [0:0] n1_idata_p0_9_;
	reg [0:0] n1_idata_p0_10_;
	reg [0:0] n1_idata_p0_11_;
	reg [0:0] n1_idata_p0_12_;
	reg [0:0] n1_idata_p0_13_;
	reg [0:0] n1_idata_p0_14_;
	reg [0:0] n1_idata_p0_15_;
	reg [0:0] n1_idata_p0_16_;
	reg [0:0] n1_idata_p0_17_;
	reg [0:0] n1_idata_p0_18_;
	reg [0:0] n1_idata_p0_19_;
	reg [0:0] n1_idata_p0_20_;
	reg [0:0] n1_idata_p0_21_;
	reg [0:0] n1_idata_p0_22_;
	reg [0:0] n1_idata_p0_23_;
	reg [0:0] n1_idata_p0_24_;
	reg [0:0] n1_idata_p0_25_;
	reg [0:0] n1_idata_p0_26_;
	reg [0:0] n1_idata_p0_27_;
	reg [0:0] n1_idata_p0_28_;
	reg [0:0] n1_idata_p0_29_;
	reg [0:0] n1_idata_p0_30_;
	reg [0:0] n1_idata_p0_31_;
	reg [0:0] n1_idata_p0_32_;
	reg [0:0] n1_idata_p0_33_;
	reg [0:0] n1_idata_p0_34_;
	reg [0:0] n1_ivalid_p0;
	reg [0:0] n1_ivch_p0;
	reg [0:0] n2_idata_p0_0_;
	reg [0:0] n2_idata_p0_1_;
	reg [0:0] n2_idata_p0_2_;
	reg [0:0] n2_idata_p0_3_;
	reg [0:0] n2_idata_p0_4_;
	reg [0:0] n2_idata_p0_5_;
	reg [0:0] n2_idata_p0_6_;
	reg [0:0] n2_idata_p0_7_;
	reg [0:0] n2_idata_p0_8_;
	reg [0:0] n2_idata_p0_9_;
	reg [0:0] n2_idata_p0_10_;
	reg [0:0] n2_idata_p0_11_;
	reg [0:0] n2_idata_p0_12_;
	reg [0:0] n2_idata_p0_13_;
	reg [0:0] n2_idata_p0_14_;
	reg [0:0] n2_idata_p0_15_;
	reg [0:0] n2_idata_p0_16_;
	reg [0:0] n2_idata_p0_17_;
	reg [0:0] n2_idata_p0_18_;
	reg [0:0] n2_idata_p0_19_;
	reg [0:0] n2_idata_p0_20_;
	reg [0:0] n2_idata_p0_21_;
	reg [0:0] n2_idata_p0_22_;
	reg [0:0] n2_idata_p0_23_;
	reg [0:0] n2_idata_p0_24_;
	reg [0:0] n2_idata_p0_25_;
	reg [0:0] n2_idata_p0_26_;
	reg [0:0] n2_idata_p0_27_;
	reg [0:0] n2_idata_p0_28_;
	reg [0:0] n2_idata_p0_29_;
	reg [0:0] n2_idata_p0_30_;
	reg [0:0] n2_idata_p0_31_;
	reg [0:0] n2_idata_p0_32_;
	reg [0:0] n2_idata_p0_33_;
	reg [0:0] n2_idata_p0_34_;
	reg [0:0] n2_ivalid_p0;
	reg [0:0] n2_ivch_p0;
	reg [0:0] n3_idata_p0_0_;
	reg [0:0] n3_idata_p0_1_;
	reg [0:0] n3_idata_p0_2_;
	reg [0:0] n3_idata_p0_3_;
	reg [0:0] n3_idata_p0_4_;
	reg [0:0] n3_idata_p0_5_;
	reg [0:0] n3_idata_p0_6_;
	reg [0:0] n3_idata_p0_7_;
	reg [0:0] n3_idata_p0_8_;
	reg [0:0] n3_idata_p0_9_;
	reg [0:0] n3_idata_p0_10_;
	reg [0:0] n3_idata_p0_11_;
	reg [0:0] n3_idata_p0_12_;
	reg [0:0] n3_idata_p0_13_;
	reg [0:0] n3_idata_p0_14_;
	reg [0:0] n3_idata_p0_15_;
	reg [0:0] n3_idata_p0_16_;
	reg [0:0] n3_idata_p0_17_;
	reg [0:0] n3_idata_p0_18_;
	reg [0:0] n3_idata_p0_19_;
	reg [0:0] n3_idata_p0_20_;
	reg [0:0] n3_idata_p0_21_;
	reg [0:0] n3_idata_p0_22_;
	reg [0:0] n3_idata_p0_23_;
	reg [0:0] n3_idata_p0_24_;
	reg [0:0] n3_idata_p0_25_;
	reg [0:0] n3_idata_p0_26_;
	reg [0:0] n3_idata_p0_27_;
	reg [0:0] n3_idata_p0_28_;
	reg [0:0] n3_idata_p0_29_;
	reg [0:0] n3_idata_p0_30_;
	reg [0:0] n3_idata_p0_31_;
	reg [0:0] n3_idata_p0_32_;
	reg [0:0] n3_idata_p0_33_;
	reg [0:0] n3_idata_p0_34_;
	reg [0:0] n3_ivalid_p0;
	reg [0:0] n3_ivch_p0;
	reg [0:0] n4_idata_p0_0_;
	reg [0:0] n4_idata_p0_1_;
	reg [0:0] n4_idata_p0_2_;
	reg [0:0] n4_idata_p0_3_;
	reg [0:0] n4_idata_p0_4_;
	reg [0:0] n4_idata_p0_5_;
	reg [0:0] n4_idata_p0_6_;
	reg [0:0] n4_idata_p0_7_;
	reg [0:0] n4_idata_p0_8_;
	reg [0:0] n4_idata_p0_9_;
	reg [0:0] n4_idata_p0_10_;
	reg [0:0] n4_idata_p0_11_;
	reg [0:0] n4_idata_p0_12_;
	reg [0:0] n4_idata_p0_13_;
	reg [0:0] n4_idata_p0_14_;
	reg [0:0] n4_idata_p0_15_;
	reg [0:0] n4_idata_p0_16_;
	reg [0:0] n4_idata_p0_17_;
	reg [0:0] n4_idata_p0_18_;
	reg [0:0] n4_idata_p0_19_;
	reg [0:0] n4_idata_p0_20_;
	reg [0:0] n4_idata_p0_21_;
	reg [0:0] n4_idata_p0_22_;
	reg [0:0] n4_idata_p0_23_;
	reg [0:0] n4_idata_p0_24_;
	reg [0:0] n4_idata_p0_25_;
	reg [0:0] n4_idata_p0_26_;
	reg [0:0] n4_idata_p0_27_;
	reg [0:0] n4_idata_p0_28_;
	reg [0:0] n4_idata_p0_29_;
	reg [0:0] n4_idata_p0_30_;
	reg [0:0] n4_idata_p0_31_;
	reg [0:0] n4_idata_p0_32_;
	reg [0:0] n4_idata_p0_33_;
	reg [0:0] n4_idata_p0_34_;
	reg [0:0] n4_ivalid_p0;
	reg [0:0] n4_ivch_p0;
	reg [0:0] n5_idata_p0_0_;
	reg [0:0] n5_idata_p0_1_;
	reg [0:0] n5_idata_p0_2_;
	reg [0:0] n5_idata_p0_3_;
	reg [0:0] n5_idata_p0_4_;
	reg [0:0] n5_idata_p0_5_;
	reg [0:0] n5_idata_p0_6_;
	reg [0:0] n5_idata_p0_7_;
	reg [0:0] n5_idata_p0_8_;
	reg [0:0] n5_idata_p0_9_;
	reg [0:0] n5_idata_p0_10_;
	reg [0:0] n5_idata_p0_11_;
	reg [0:0] n5_idata_p0_12_;
	reg [0:0] n5_idata_p0_13_;
	reg [0:0] n5_idata_p0_14_;
	reg [0:0] n5_idata_p0_15_;
	reg [0:0] n5_idata_p0_16_;
	reg [0:0] n5_idata_p0_17_;
	reg [0:0] n5_idata_p0_18_;
	reg [0:0] n5_idata_p0_19_;
	reg [0:0] n5_idata_p0_20_;
	reg [0:0] n5_idata_p0_21_;
	reg [0:0] n5_idata_p0_22_;
	reg [0:0] n5_idata_p0_23_;
	reg [0:0] n5_idata_p0_24_;
	reg [0:0] n5_idata_p0_25_;
	reg [0:0] n5_idata_p0_26_;
	reg [0:0] n5_idata_p0_27_;
	reg [0:0] n5_idata_p0_28_;
	reg [0:0] n5_idata_p0_29_;
	reg [0:0] n5_idata_p0_30_;
	reg [0:0] n5_idata_p0_31_;
	reg [0:0] n5_idata_p0_32_;
	reg [0:0] n5_idata_p0_33_;
	reg [0:0] n5_idata_p0_34_;
	reg [0:0] n5_ivalid_p0;
	reg [0:0] n5_ivch_p0;
	reg [0:0] n6_idata_p0_0_;
	reg [0:0] n6_idata_p0_1_;
	reg [0:0] n6_idata_p0_2_;
	reg [0:0] n6_idata_p0_3_;
	reg [0:0] n6_idata_p0_4_;
	reg [0:0] n6_idata_p0_5_;
	reg [0:0] n6_idata_p0_6_;
	reg [0:0] n6_idata_p0_7_;
	reg [0:0] n6_idata_p0_8_;
	reg [0:0] n6_idata_p0_9_;
	reg [0:0] n6_idata_p0_10_;
	reg [0:0] n6_idata_p0_11_;
	reg [0:0] n6_idata_p0_12_;
	reg [0:0] n6_idata_p0_13_;
	reg [0:0] n6_idata_p0_14_;
	reg [0:0] n6_idata_p0_15_;
	reg [0:0] n6_idata_p0_16_;
	reg [0:0] n6_idata_p0_17_;
	reg [0:0] n6_idata_p0_18_;
	reg [0:0] n6_idata_p0_19_;
	reg [0:0] n6_idata_p0_20_;
	reg [0:0] n6_idata_p0_21_;
	reg [0:0] n6_idata_p0_22_;
	reg [0:0] n6_idata_p0_23_;
	reg [0:0] n6_idata_p0_24_;
	reg [0:0] n6_idata_p0_25_;
	reg [0:0] n6_idata_p0_26_;
	reg [0:0] n6_idata_p0_27_;
	reg [0:0] n6_idata_p0_28_;
	reg [0:0] n6_idata_p0_29_;
	reg [0:0] n6_idata_p0_30_;
	reg [0:0] n6_idata_p0_31_;
	reg [0:0] n6_idata_p0_32_;
	reg [0:0] n6_idata_p0_33_;
	reg [0:0] n6_idata_p0_34_;
	reg [0:0] n6_ivalid_p0;
	reg [0:0] n6_ivch_p0;
	reg [0:0] n7_idata_p0_0_;
	reg [0:0] n7_idata_p0_1_;
	reg [0:0] n7_idata_p0_2_;
	reg [0:0] n7_idata_p0_3_;
	reg [0:0] n7_idata_p0_4_;
	reg [0:0] n7_idata_p0_5_;
	reg [0:0] n7_idata_p0_6_;
	reg [0:0] n7_idata_p0_7_;
	reg [0:0] n7_idata_p0_8_;
	reg [0:0] n7_idata_p0_9_;
	reg [0:0] n7_idata_p0_10_;
	reg [0:0] n7_idata_p0_11_;
	reg [0:0] n7_idata_p0_12_;
	reg [0:0] n7_idata_p0_13_;
	reg [0:0] n7_idata_p0_14_;
	reg [0:0] n7_idata_p0_15_;
	reg [0:0] n7_idata_p0_16_;
	reg [0:0] n7_idata_p0_17_;
	reg [0:0] n7_idata_p0_18_;
	reg [0:0] n7_idata_p0_19_;
	reg [0:0] n7_idata_p0_20_;
	reg [0:0] n7_idata_p0_21_;
	reg [0:0] n7_idata_p0_22_;
	reg [0:0] n7_idata_p0_23_;
	reg [0:0] n7_idata_p0_24_;
	reg [0:0] n7_idata_p0_25_;
	reg [0:0] n7_idata_p0_26_;
	reg [0:0] n7_idata_p0_27_;
	reg [0:0] n7_idata_p0_28_;
	reg [0:0] n7_idata_p0_29_;
	reg [0:0] n7_idata_p0_30_;
	reg [0:0] n7_idata_p0_31_;
	reg [0:0] n7_idata_p0_32_;
	reg [0:0] n7_idata_p0_33_;
	reg [0:0] n7_idata_p0_34_;
	reg [0:0] n7_ivalid_p0;
	reg [0:0] n7_ivch_p0;
	reg [0:0] n8_idata_p0_0_;
	reg [0:0] n8_idata_p0_1_;
	reg [0:0] n8_idata_p0_2_;
	reg [0:0] n8_idata_p0_3_;
	reg [0:0] n8_idata_p0_4_;
	reg [0:0] n8_idata_p0_5_;
	reg [0:0] n8_idata_p0_6_;
	reg [0:0] n8_idata_p0_7_;
	reg [0:0] n8_idata_p0_8_;
	reg [0:0] n8_idata_p0_9_;
	reg [0:0] n8_idata_p0_10_;
	reg [0:0] n8_idata_p0_11_;
	reg [0:0] n8_idata_p0_12_;
	reg [0:0] n8_idata_p0_13_;
	reg [0:0] n8_idata_p0_14_;
	reg [0:0] n8_idata_p0_15_;
	reg [0:0] n8_idata_p0_16_;
	reg [0:0] n8_idata_p0_17_;
	reg [0:0] n8_idata_p0_18_;
	reg [0:0] n8_idata_p0_19_;
	reg [0:0] n8_idata_p0_20_;
	reg [0:0] n8_idata_p0_21_;
	reg [0:0] n8_idata_p0_22_;
	reg [0:0] n8_idata_p0_23_;
	reg [0:0] n8_idata_p0_24_;
	reg [0:0] n8_idata_p0_25_;
	reg [0:0] n8_idata_p0_26_;
	reg [0:0] n8_idata_p0_27_;
	reg [0:0] n8_idata_p0_28_;
	reg [0:0] n8_idata_p0_29_;
	reg [0:0] n8_idata_p0_30_;
	reg [0:0] n8_idata_p0_31_;
	reg [0:0] n8_idata_p0_32_;
	reg [0:0] n8_idata_p0_33_;
	reg [0:0] n8_idata_p0_34_;
	reg [0:0] n8_ivalid_p0;
	reg [0:0] n8_ivch_p0;
	reg [0:0] rst_;

// ----- FPGA fabric outputs -------
	wire [0:0] n0_ordy_p0_0__gfpga;
	wire [0:0] n0_ordy_p0_1__gfpga;
	wire [0:0] n0_odata_p0_0__gfpga;
	wire [0:0] n0_odata_p0_1__gfpga;
	wire [0:0] n0_odata_p0_2__gfpga;
	wire [0:0] n0_odata_p0_3__gfpga;
	wire [0:0] n0_odata_p0_4__gfpga;
	wire [0:0] n0_odata_p0_5__gfpga;
	wire [0:0] n0_odata_p0_6__gfpga;
	wire [0:0] n0_odata_p0_7__gfpga;
	wire [0:0] n0_odata_p0_8__gfpga;
	wire [0:0] n0_odata_p0_9__gfpga;
	wire [0:0] n0_odata_p0_10__gfpga;
	wire [0:0] n0_odata_p0_11__gfpga;
	wire [0:0] n0_odata_p0_12__gfpga;
	wire [0:0] n0_odata_p0_13__gfpga;
	wire [0:0] n0_odata_p0_14__gfpga;
	wire [0:0] n0_odata_p0_15__gfpga;
	wire [0:0] n0_odata_p0_16__gfpga;
	wire [0:0] n0_odata_p0_17__gfpga;
	wire [0:0] n0_odata_p0_18__gfpga;
	wire [0:0] n0_odata_p0_19__gfpga;
	wire [0:0] n0_odata_p0_20__gfpga;
	wire [0:0] n0_odata_p0_21__gfpga;
	wire [0:0] n0_odata_p0_22__gfpga;
	wire [0:0] n0_odata_p0_23__gfpga;
	wire [0:0] n0_odata_p0_24__gfpga;
	wire [0:0] n0_odata_p0_25__gfpga;
	wire [0:0] n0_odata_p0_26__gfpga;
	wire [0:0] n0_odata_p0_27__gfpga;
	wire [0:0] n0_odata_p0_28__gfpga;
	wire [0:0] n0_odata_p0_29__gfpga;
	wire [0:0] n0_odata_p0_30__gfpga;
	wire [0:0] n0_odata_p0_31__gfpga;
	wire [0:0] n0_odata_p0_32__gfpga;
	wire [0:0] n0_odata_p0_33__gfpga;
	wire [0:0] n0_odata_p0_34__gfpga;
	wire [0:0] n0_ovalid_p0_gfpga;
	wire [0:0] n1_ordy_p0_0__gfpga;
	wire [0:0] n1_ordy_p0_1__gfpga;
	wire [0:0] n1_odata_p0_0__gfpga;
	wire [0:0] n1_odata_p0_1__gfpga;
	wire [0:0] n1_odata_p0_2__gfpga;
	wire [0:0] n1_odata_p0_3__gfpga;
	wire [0:0] n1_odata_p0_4__gfpga;
	wire [0:0] n1_odata_p0_5__gfpga;
	wire [0:0] n1_odata_p0_6__gfpga;
	wire [0:0] n1_odata_p0_7__gfpga;
	wire [0:0] n1_odata_p0_8__gfpga;
	wire [0:0] n1_odata_p0_9__gfpga;
	wire [0:0] n1_odata_p0_10__gfpga;
	wire [0:0] n1_odata_p0_11__gfpga;
	wire [0:0] n1_odata_p0_12__gfpga;
	wire [0:0] n1_odata_p0_13__gfpga;
	wire [0:0] n1_odata_p0_14__gfpga;
	wire [0:0] n1_odata_p0_15__gfpga;
	wire [0:0] n1_odata_p0_16__gfpga;
	wire [0:0] n1_odata_p0_17__gfpga;
	wire [0:0] n1_odata_p0_18__gfpga;
	wire [0:0] n1_odata_p0_19__gfpga;
	wire [0:0] n1_odata_p0_20__gfpga;
	wire [0:0] n1_odata_p0_21__gfpga;
	wire [0:0] n1_odata_p0_22__gfpga;
	wire [0:0] n1_odata_p0_23__gfpga;
	wire [0:0] n1_odata_p0_24__gfpga;
	wire [0:0] n1_odata_p0_25__gfpga;
	wire [0:0] n1_odata_p0_26__gfpga;
	wire [0:0] n1_odata_p0_27__gfpga;
	wire [0:0] n1_odata_p0_28__gfpga;
	wire [0:0] n1_odata_p0_29__gfpga;
	wire [0:0] n1_odata_p0_30__gfpga;
	wire [0:0] n1_odata_p0_31__gfpga;
	wire [0:0] n1_odata_p0_32__gfpga;
	wire [0:0] n1_odata_p0_33__gfpga;
	wire [0:0] n1_odata_p0_34__gfpga;
	wire [0:0] n1_ovalid_p0_gfpga;
	wire [0:0] n2_ordy_p0_0__gfpga;
	wire [0:0] n2_ordy_p0_1__gfpga;
	wire [0:0] n2_odata_p0_0__gfpga;
	wire [0:0] n2_odata_p0_1__gfpga;
	wire [0:0] n2_odata_p0_2__gfpga;
	wire [0:0] n2_odata_p0_3__gfpga;
	wire [0:0] n2_odata_p0_4__gfpga;
	wire [0:0] n2_odata_p0_5__gfpga;
	wire [0:0] n2_odata_p0_6__gfpga;
	wire [0:0] n2_odata_p0_7__gfpga;
	wire [0:0] n2_odata_p0_8__gfpga;
	wire [0:0] n2_odata_p0_9__gfpga;
	wire [0:0] n2_odata_p0_10__gfpga;
	wire [0:0] n2_odata_p0_11__gfpga;
	wire [0:0] n2_odata_p0_12__gfpga;
	wire [0:0] n2_odata_p0_13__gfpga;
	wire [0:0] n2_odata_p0_14__gfpga;
	wire [0:0] n2_odata_p0_15__gfpga;
	wire [0:0] n2_odata_p0_16__gfpga;
	wire [0:0] n2_odata_p0_17__gfpga;
	wire [0:0] n2_odata_p0_18__gfpga;
	wire [0:0] n2_odata_p0_19__gfpga;
	wire [0:0] n2_odata_p0_20__gfpga;
	wire [0:0] n2_odata_p0_21__gfpga;
	wire [0:0] n2_odata_p0_22__gfpga;
	wire [0:0] n2_odata_p0_23__gfpga;
	wire [0:0] n2_odata_p0_24__gfpga;
	wire [0:0] n2_odata_p0_25__gfpga;
	wire [0:0] n2_odata_p0_26__gfpga;
	wire [0:0] n2_odata_p0_27__gfpga;
	wire [0:0] n2_odata_p0_28__gfpga;
	wire [0:0] n2_odata_p0_29__gfpga;
	wire [0:0] n2_odata_p0_30__gfpga;
	wire [0:0] n2_odata_p0_31__gfpga;
	wire [0:0] n2_odata_p0_32__gfpga;
	wire [0:0] n2_odata_p0_33__gfpga;
	wire [0:0] n2_odata_p0_34__gfpga;
	wire [0:0] n2_ovalid_p0_gfpga;
	wire [0:0] n3_ordy_p0_0__gfpga;
	wire [0:0] n3_ordy_p0_1__gfpga;
	wire [0:0] n3_odata_p0_0__gfpga;
	wire [0:0] n3_odata_p0_1__gfpga;
	wire [0:0] n3_odata_p0_2__gfpga;
	wire [0:0] n3_odata_p0_3__gfpga;
	wire [0:0] n3_odata_p0_4__gfpga;
	wire [0:0] n3_odata_p0_5__gfpga;
	wire [0:0] n3_odata_p0_6__gfpga;
	wire [0:0] n3_odata_p0_7__gfpga;
	wire [0:0] n3_odata_p0_8__gfpga;
	wire [0:0] n3_odata_p0_9__gfpga;
	wire [0:0] n3_odata_p0_10__gfpga;
	wire [0:0] n3_odata_p0_11__gfpga;
	wire [0:0] n3_odata_p0_12__gfpga;
	wire [0:0] n3_odata_p0_13__gfpga;
	wire [0:0] n3_odata_p0_14__gfpga;
	wire [0:0] n3_odata_p0_15__gfpga;
	wire [0:0] n3_odata_p0_16__gfpga;
	wire [0:0] n3_odata_p0_17__gfpga;
	wire [0:0] n3_odata_p0_18__gfpga;
	wire [0:0] n3_odata_p0_19__gfpga;
	wire [0:0] n3_odata_p0_20__gfpga;
	wire [0:0] n3_odata_p0_21__gfpga;
	wire [0:0] n3_odata_p0_22__gfpga;
	wire [0:0] n3_odata_p0_23__gfpga;
	wire [0:0] n3_odata_p0_24__gfpga;
	wire [0:0] n3_odata_p0_25__gfpga;
	wire [0:0] n3_odata_p0_26__gfpga;
	wire [0:0] n3_odata_p0_27__gfpga;
	wire [0:0] n3_odata_p0_28__gfpga;
	wire [0:0] n3_odata_p0_29__gfpga;
	wire [0:0] n3_odata_p0_30__gfpga;
	wire [0:0] n3_odata_p0_31__gfpga;
	wire [0:0] n3_odata_p0_32__gfpga;
	wire [0:0] n3_odata_p0_33__gfpga;
	wire [0:0] n3_odata_p0_34__gfpga;
	wire [0:0] n3_ovalid_p0_gfpga;
	wire [0:0] n4_ordy_p0_0__gfpga;
	wire [0:0] n4_ordy_p0_1__gfpga;
	wire [0:0] n4_odata_p0_0__gfpga;
	wire [0:0] n4_odata_p0_1__gfpga;
	wire [0:0] n4_odata_p0_2__gfpga;
	wire [0:0] n4_odata_p0_3__gfpga;
	wire [0:0] n4_odata_p0_4__gfpga;
	wire [0:0] n4_odata_p0_5__gfpga;
	wire [0:0] n4_odata_p0_6__gfpga;
	wire [0:0] n4_odata_p0_7__gfpga;
	wire [0:0] n4_odata_p0_8__gfpga;
	wire [0:0] n4_odata_p0_9__gfpga;
	wire [0:0] n4_odata_p0_10__gfpga;
	wire [0:0] n4_odata_p0_11__gfpga;
	wire [0:0] n4_odata_p0_12__gfpga;
	wire [0:0] n4_odata_p0_13__gfpga;
	wire [0:0] n4_odata_p0_14__gfpga;
	wire [0:0] n4_odata_p0_15__gfpga;
	wire [0:0] n4_odata_p0_16__gfpga;
	wire [0:0] n4_odata_p0_17__gfpga;
	wire [0:0] n4_odata_p0_18__gfpga;
	wire [0:0] n4_odata_p0_19__gfpga;
	wire [0:0] n4_odata_p0_20__gfpga;
	wire [0:0] n4_odata_p0_21__gfpga;
	wire [0:0] n4_odata_p0_22__gfpga;
	wire [0:0] n4_odata_p0_23__gfpga;
	wire [0:0] n4_odata_p0_24__gfpga;
	wire [0:0] n4_odata_p0_25__gfpga;
	wire [0:0] n4_odata_p0_26__gfpga;
	wire [0:0] n4_odata_p0_27__gfpga;
	wire [0:0] n4_odata_p0_28__gfpga;
	wire [0:0] n4_odata_p0_29__gfpga;
	wire [0:0] n4_odata_p0_30__gfpga;
	wire [0:0] n4_odata_p0_31__gfpga;
	wire [0:0] n4_odata_p0_32__gfpga;
	wire [0:0] n4_odata_p0_33__gfpga;
	wire [0:0] n4_odata_p0_34__gfpga;
	wire [0:0] n4_ovalid_p0_gfpga;
	wire [0:0] n5_ordy_p0_0__gfpga;
	wire [0:0] n5_ordy_p0_1__gfpga;
	wire [0:0] n5_odata_p0_0__gfpga;
	wire [0:0] n5_odata_p0_1__gfpga;
	wire [0:0] n5_odata_p0_2__gfpga;
	wire [0:0] n5_odata_p0_3__gfpga;
	wire [0:0] n5_odata_p0_4__gfpga;
	wire [0:0] n5_odata_p0_5__gfpga;
	wire [0:0] n5_odata_p0_6__gfpga;
	wire [0:0] n5_odata_p0_7__gfpga;
	wire [0:0] n5_odata_p0_8__gfpga;
	wire [0:0] n5_odata_p0_9__gfpga;
	wire [0:0] n5_odata_p0_10__gfpga;
	wire [0:0] n5_odata_p0_11__gfpga;
	wire [0:0] n5_odata_p0_12__gfpga;
	wire [0:0] n5_odata_p0_13__gfpga;
	wire [0:0] n5_odata_p0_14__gfpga;
	wire [0:0] n5_odata_p0_15__gfpga;
	wire [0:0] n5_odata_p0_16__gfpga;
	wire [0:0] n5_odata_p0_17__gfpga;
	wire [0:0] n5_odata_p0_18__gfpga;
	wire [0:0] n5_odata_p0_19__gfpga;
	wire [0:0] n5_odata_p0_20__gfpga;
	wire [0:0] n5_odata_p0_21__gfpga;
	wire [0:0] n5_odata_p0_22__gfpga;
	wire [0:0] n5_odata_p0_23__gfpga;
	wire [0:0] n5_odata_p0_24__gfpga;
	wire [0:0] n5_odata_p0_25__gfpga;
	wire [0:0] n5_odata_p0_26__gfpga;
	wire [0:0] n5_odata_p0_27__gfpga;
	wire [0:0] n5_odata_p0_28__gfpga;
	wire [0:0] n5_odata_p0_29__gfpga;
	wire [0:0] n5_odata_p0_30__gfpga;
	wire [0:0] n5_odata_p0_31__gfpga;
	wire [0:0] n5_odata_p0_32__gfpga;
	wire [0:0] n5_odata_p0_33__gfpga;
	wire [0:0] n5_odata_p0_34__gfpga;
	wire [0:0] n5_ovalid_p0_gfpga;
	wire [0:0] n6_ordy_p0_0__gfpga;
	wire [0:0] n6_ordy_p0_1__gfpga;
	wire [0:0] n6_odata_p0_0__gfpga;
	wire [0:0] n6_odata_p0_1__gfpga;
	wire [0:0] n6_odata_p0_2__gfpga;
	wire [0:0] n6_odata_p0_3__gfpga;
	wire [0:0] n6_odata_p0_4__gfpga;
	wire [0:0] n6_odata_p0_5__gfpga;
	wire [0:0] n6_odata_p0_6__gfpga;
	wire [0:0] n6_odata_p0_7__gfpga;
	wire [0:0] n6_odata_p0_8__gfpga;
	wire [0:0] n6_odata_p0_9__gfpga;
	wire [0:0] n6_odata_p0_10__gfpga;
	wire [0:0] n6_odata_p0_11__gfpga;
	wire [0:0] n6_odata_p0_12__gfpga;
	wire [0:0] n6_odata_p0_13__gfpga;
	wire [0:0] n6_odata_p0_14__gfpga;
	wire [0:0] n6_odata_p0_15__gfpga;
	wire [0:0] n6_odata_p0_16__gfpga;
	wire [0:0] n6_odata_p0_17__gfpga;
	wire [0:0] n6_odata_p0_18__gfpga;
	wire [0:0] n6_odata_p0_19__gfpga;
	wire [0:0] n6_odata_p0_20__gfpga;
	wire [0:0] n6_odata_p0_21__gfpga;
	wire [0:0] n6_odata_p0_22__gfpga;
	wire [0:0] n6_odata_p0_23__gfpga;
	wire [0:0] n6_odata_p0_24__gfpga;
	wire [0:0] n6_odata_p0_25__gfpga;
	wire [0:0] n6_odata_p0_26__gfpga;
	wire [0:0] n6_odata_p0_27__gfpga;
	wire [0:0] n6_odata_p0_28__gfpga;
	wire [0:0] n6_odata_p0_29__gfpga;
	wire [0:0] n6_odata_p0_30__gfpga;
	wire [0:0] n6_odata_p0_31__gfpga;
	wire [0:0] n6_odata_p0_32__gfpga;
	wire [0:0] n6_odata_p0_33__gfpga;
	wire [0:0] n6_odata_p0_34__gfpga;
	wire [0:0] n6_ovalid_p0_gfpga;
	wire [0:0] n7_ordy_p0_0__gfpga;
	wire [0:0] n7_ordy_p0_1__gfpga;
	wire [0:0] n7_odata_p0_0__gfpga;
	wire [0:0] n7_odata_p0_1__gfpga;
	wire [0:0] n7_odata_p0_2__gfpga;
	wire [0:0] n7_odata_p0_3__gfpga;
	wire [0:0] n7_odata_p0_4__gfpga;
	wire [0:0] n7_odata_p0_5__gfpga;
	wire [0:0] n7_odata_p0_6__gfpga;
	wire [0:0] n7_odata_p0_7__gfpga;
	wire [0:0] n7_odata_p0_8__gfpga;
	wire [0:0] n7_odata_p0_9__gfpga;
	wire [0:0] n7_odata_p0_10__gfpga;
	wire [0:0] n7_odata_p0_11__gfpga;
	wire [0:0] n7_odata_p0_12__gfpga;
	wire [0:0] n7_odata_p0_13__gfpga;
	wire [0:0] n7_odata_p0_14__gfpga;
	wire [0:0] n7_odata_p0_15__gfpga;
	wire [0:0] n7_odata_p0_16__gfpga;
	wire [0:0] n7_odata_p0_17__gfpga;
	wire [0:0] n7_odata_p0_18__gfpga;
	wire [0:0] n7_odata_p0_19__gfpga;
	wire [0:0] n7_odata_p0_20__gfpga;
	wire [0:0] n7_odata_p0_21__gfpga;
	wire [0:0] n7_odata_p0_22__gfpga;
	wire [0:0] n7_odata_p0_23__gfpga;
	wire [0:0] n7_odata_p0_24__gfpga;
	wire [0:0] n7_odata_p0_25__gfpga;
	wire [0:0] n7_odata_p0_26__gfpga;
	wire [0:0] n7_odata_p0_27__gfpga;
	wire [0:0] n7_odata_p0_28__gfpga;
	wire [0:0] n7_odata_p0_29__gfpga;
	wire [0:0] n7_odata_p0_30__gfpga;
	wire [0:0] n7_odata_p0_31__gfpga;
	wire [0:0] n7_odata_p0_32__gfpga;
	wire [0:0] n7_odata_p0_33__gfpga;
	wire [0:0] n7_odata_p0_34__gfpga;
	wire [0:0] n7_ovalid_p0_gfpga;
	wire [0:0] n8_ordy_p0_0__gfpga;
	wire [0:0] n8_ordy_p0_1__gfpga;
	wire [0:0] n8_odata_p0_0__gfpga;
	wire [0:0] n8_odata_p0_1__gfpga;
	wire [0:0] n8_odata_p0_2__gfpga;
	wire [0:0] n8_odata_p0_3__gfpga;
	wire [0:0] n8_odata_p0_4__gfpga;
	wire [0:0] n8_odata_p0_5__gfpga;
	wire [0:0] n8_odata_p0_6__gfpga;
	wire [0:0] n8_odata_p0_7__gfpga;
	wire [0:0] n8_odata_p0_8__gfpga;
	wire [0:0] n8_odata_p0_9__gfpga;
	wire [0:0] n8_odata_p0_10__gfpga;
	wire [0:0] n8_odata_p0_11__gfpga;
	wire [0:0] n8_odata_p0_12__gfpga;
	wire [0:0] n8_odata_p0_13__gfpga;
	wire [0:0] n8_odata_p0_14__gfpga;
	wire [0:0] n8_odata_p0_15__gfpga;
	wire [0:0] n8_odata_p0_16__gfpga;
	wire [0:0] n8_odata_p0_17__gfpga;
	wire [0:0] n8_odata_p0_18__gfpga;
	wire [0:0] n8_odata_p0_19__gfpga;
	wire [0:0] n8_odata_p0_20__gfpga;
	wire [0:0] n8_odata_p0_21__gfpga;
	wire [0:0] n8_odata_p0_22__gfpga;
	wire [0:0] n8_odata_p0_23__gfpga;
	wire [0:0] n8_odata_p0_24__gfpga;
	wire [0:0] n8_odata_p0_25__gfpga;
	wire [0:0] n8_odata_p0_26__gfpga;
	wire [0:0] n8_odata_p0_27__gfpga;
	wire [0:0] n8_odata_p0_28__gfpga;
	wire [0:0] n8_odata_p0_29__gfpga;
	wire [0:0] n8_odata_p0_30__gfpga;
	wire [0:0] n8_odata_p0_31__gfpga;
	wire [0:0] n8_odata_p0_32__gfpga;
	wire [0:0] n8_odata_p0_33__gfpga;
	wire [0:0] n8_odata_p0_34__gfpga;
	wire [0:0] n8_ovalid_p0_gfpga;

// ----- Benchmark outputs -------
	wire [0:0] n0_ordy_p0_0__bench;
	wire [0:0] n0_ordy_p0_1__bench;
	wire [0:0] n0_odata_p0_0__bench;
	wire [0:0] n0_odata_p0_1__bench;
	wire [0:0] n0_odata_p0_2__bench;
	wire [0:0] n0_odata_p0_3__bench;
	wire [0:0] n0_odata_p0_4__bench;
	wire [0:0] n0_odata_p0_5__bench;
	wire [0:0] n0_odata_p0_6__bench;
	wire [0:0] n0_odata_p0_7__bench;
	wire [0:0] n0_odata_p0_8__bench;
	wire [0:0] n0_odata_p0_9__bench;
	wire [0:0] n0_odata_p0_10__bench;
	wire [0:0] n0_odata_p0_11__bench;
	wire [0:0] n0_odata_p0_12__bench;
	wire [0:0] n0_odata_p0_13__bench;
	wire [0:0] n0_odata_p0_14__bench;
	wire [0:0] n0_odata_p0_15__bench;
	wire [0:0] n0_odata_p0_16__bench;
	wire [0:0] n0_odata_p0_17__bench;
	wire [0:0] n0_odata_p0_18__bench;
	wire [0:0] n0_odata_p0_19__bench;
	wire [0:0] n0_odata_p0_20__bench;
	wire [0:0] n0_odata_p0_21__bench;
	wire [0:0] n0_odata_p0_22__bench;
	wire [0:0] n0_odata_p0_23__bench;
	wire [0:0] n0_odata_p0_24__bench;
	wire [0:0] n0_odata_p0_25__bench;
	wire [0:0] n0_odata_p0_26__bench;
	wire [0:0] n0_odata_p0_27__bench;
	wire [0:0] n0_odata_p0_28__bench;
	wire [0:0] n0_odata_p0_29__bench;
	wire [0:0] n0_odata_p0_30__bench;
	wire [0:0] n0_odata_p0_31__bench;
	wire [0:0] n0_odata_p0_32__bench;
	wire [0:0] n0_odata_p0_33__bench;
	wire [0:0] n0_odata_p0_34__bench;
	wire [0:0] n0_ovalid_p0_bench;
	wire [0:0] n1_ordy_p0_0__bench;
	wire [0:0] n1_ordy_p0_1__bench;
	wire [0:0] n1_odata_p0_0__bench;
	wire [0:0] n1_odata_p0_1__bench;
	wire [0:0] n1_odata_p0_2__bench;
	wire [0:0] n1_odata_p0_3__bench;
	wire [0:0] n1_odata_p0_4__bench;
	wire [0:0] n1_odata_p0_5__bench;
	wire [0:0] n1_odata_p0_6__bench;
	wire [0:0] n1_odata_p0_7__bench;
	wire [0:0] n1_odata_p0_8__bench;
	wire [0:0] n1_odata_p0_9__bench;
	wire [0:0] n1_odata_p0_10__bench;
	wire [0:0] n1_odata_p0_11__bench;
	wire [0:0] n1_odata_p0_12__bench;
	wire [0:0] n1_odata_p0_13__bench;
	wire [0:0] n1_odata_p0_14__bench;
	wire [0:0] n1_odata_p0_15__bench;
	wire [0:0] n1_odata_p0_16__bench;
	wire [0:0] n1_odata_p0_17__bench;
	wire [0:0] n1_odata_p0_18__bench;
	wire [0:0] n1_odata_p0_19__bench;
	wire [0:0] n1_odata_p0_20__bench;
	wire [0:0] n1_odata_p0_21__bench;
	wire [0:0] n1_odata_p0_22__bench;
	wire [0:0] n1_odata_p0_23__bench;
	wire [0:0] n1_odata_p0_24__bench;
	wire [0:0] n1_odata_p0_25__bench;
	wire [0:0] n1_odata_p0_26__bench;
	wire [0:0] n1_odata_p0_27__bench;
	wire [0:0] n1_odata_p0_28__bench;
	wire [0:0] n1_odata_p0_29__bench;
	wire [0:0] n1_odata_p0_30__bench;
	wire [0:0] n1_odata_p0_31__bench;
	wire [0:0] n1_odata_p0_32__bench;
	wire [0:0] n1_odata_p0_33__bench;
	wire [0:0] n1_odata_p0_34__bench;
	wire [0:0] n1_ovalid_p0_bench;
	wire [0:0] n2_ordy_p0_0__bench;
	wire [0:0] n2_ordy_p0_1__bench;
	wire [0:0] n2_odata_p0_0__bench;
	wire [0:0] n2_odata_p0_1__bench;
	wire [0:0] n2_odata_p0_2__bench;
	wire [0:0] n2_odata_p0_3__bench;
	wire [0:0] n2_odata_p0_4__bench;
	wire [0:0] n2_odata_p0_5__bench;
	wire [0:0] n2_odata_p0_6__bench;
	wire [0:0] n2_odata_p0_7__bench;
	wire [0:0] n2_odata_p0_8__bench;
	wire [0:0] n2_odata_p0_9__bench;
	wire [0:0] n2_odata_p0_10__bench;
	wire [0:0] n2_odata_p0_11__bench;
	wire [0:0] n2_odata_p0_12__bench;
	wire [0:0] n2_odata_p0_13__bench;
	wire [0:0] n2_odata_p0_14__bench;
	wire [0:0] n2_odata_p0_15__bench;
	wire [0:0] n2_odata_p0_16__bench;
	wire [0:0] n2_odata_p0_17__bench;
	wire [0:0] n2_odata_p0_18__bench;
	wire [0:0] n2_odata_p0_19__bench;
	wire [0:0] n2_odata_p0_20__bench;
	wire [0:0] n2_odata_p0_21__bench;
	wire [0:0] n2_odata_p0_22__bench;
	wire [0:0] n2_odata_p0_23__bench;
	wire [0:0] n2_odata_p0_24__bench;
	wire [0:0] n2_odata_p0_25__bench;
	wire [0:0] n2_odata_p0_26__bench;
	wire [0:0] n2_odata_p0_27__bench;
	wire [0:0] n2_odata_p0_28__bench;
	wire [0:0] n2_odata_p0_29__bench;
	wire [0:0] n2_odata_p0_30__bench;
	wire [0:0] n2_odata_p0_31__bench;
	wire [0:0] n2_odata_p0_32__bench;
	wire [0:0] n2_odata_p0_33__bench;
	wire [0:0] n2_odata_p0_34__bench;
	wire [0:0] n2_ovalid_p0_bench;
	wire [0:0] n3_ordy_p0_0__bench;
	wire [0:0] n3_ordy_p0_1__bench;
	wire [0:0] n3_odata_p0_0__bench;
	wire [0:0] n3_odata_p0_1__bench;
	wire [0:0] n3_odata_p0_2__bench;
	wire [0:0] n3_odata_p0_3__bench;
	wire [0:0] n3_odata_p0_4__bench;
	wire [0:0] n3_odata_p0_5__bench;
	wire [0:0] n3_odata_p0_6__bench;
	wire [0:0] n3_odata_p0_7__bench;
	wire [0:0] n3_odata_p0_8__bench;
	wire [0:0] n3_odata_p0_9__bench;
	wire [0:0] n3_odata_p0_10__bench;
	wire [0:0] n3_odata_p0_11__bench;
	wire [0:0] n3_odata_p0_12__bench;
	wire [0:0] n3_odata_p0_13__bench;
	wire [0:0] n3_odata_p0_14__bench;
	wire [0:0] n3_odata_p0_15__bench;
	wire [0:0] n3_odata_p0_16__bench;
	wire [0:0] n3_odata_p0_17__bench;
	wire [0:0] n3_odata_p0_18__bench;
	wire [0:0] n3_odata_p0_19__bench;
	wire [0:0] n3_odata_p0_20__bench;
	wire [0:0] n3_odata_p0_21__bench;
	wire [0:0] n3_odata_p0_22__bench;
	wire [0:0] n3_odata_p0_23__bench;
	wire [0:0] n3_odata_p0_24__bench;
	wire [0:0] n3_odata_p0_25__bench;
	wire [0:0] n3_odata_p0_26__bench;
	wire [0:0] n3_odata_p0_27__bench;
	wire [0:0] n3_odata_p0_28__bench;
	wire [0:0] n3_odata_p0_29__bench;
	wire [0:0] n3_odata_p0_30__bench;
	wire [0:0] n3_odata_p0_31__bench;
	wire [0:0] n3_odata_p0_32__bench;
	wire [0:0] n3_odata_p0_33__bench;
	wire [0:0] n3_odata_p0_34__bench;
	wire [0:0] n3_ovalid_p0_bench;
	wire [0:0] n4_ordy_p0_0__bench;
	wire [0:0] n4_ordy_p0_1__bench;
	wire [0:0] n4_odata_p0_0__bench;
	wire [0:0] n4_odata_p0_1__bench;
	wire [0:0] n4_odata_p0_2__bench;
	wire [0:0] n4_odata_p0_3__bench;
	wire [0:0] n4_odata_p0_4__bench;
	wire [0:0] n4_odata_p0_5__bench;
	wire [0:0] n4_odata_p0_6__bench;
	wire [0:0] n4_odata_p0_7__bench;
	wire [0:0] n4_odata_p0_8__bench;
	wire [0:0] n4_odata_p0_9__bench;
	wire [0:0] n4_odata_p0_10__bench;
	wire [0:0] n4_odata_p0_11__bench;
	wire [0:0] n4_odata_p0_12__bench;
	wire [0:0] n4_odata_p0_13__bench;
	wire [0:0] n4_odata_p0_14__bench;
	wire [0:0] n4_odata_p0_15__bench;
	wire [0:0] n4_odata_p0_16__bench;
	wire [0:0] n4_odata_p0_17__bench;
	wire [0:0] n4_odata_p0_18__bench;
	wire [0:0] n4_odata_p0_19__bench;
	wire [0:0] n4_odata_p0_20__bench;
	wire [0:0] n4_odata_p0_21__bench;
	wire [0:0] n4_odata_p0_22__bench;
	wire [0:0] n4_odata_p0_23__bench;
	wire [0:0] n4_odata_p0_24__bench;
	wire [0:0] n4_odata_p0_25__bench;
	wire [0:0] n4_odata_p0_26__bench;
	wire [0:0] n4_odata_p0_27__bench;
	wire [0:0] n4_odata_p0_28__bench;
	wire [0:0] n4_odata_p0_29__bench;
	wire [0:0] n4_odata_p0_30__bench;
	wire [0:0] n4_odata_p0_31__bench;
	wire [0:0] n4_odata_p0_32__bench;
	wire [0:0] n4_odata_p0_33__bench;
	wire [0:0] n4_odata_p0_34__bench;
	wire [0:0] n4_ovalid_p0_bench;
	wire [0:0] n5_ordy_p0_0__bench;
	wire [0:0] n5_ordy_p0_1__bench;
	wire [0:0] n5_odata_p0_0__bench;
	wire [0:0] n5_odata_p0_1__bench;
	wire [0:0] n5_odata_p0_2__bench;
	wire [0:0] n5_odata_p0_3__bench;
	wire [0:0] n5_odata_p0_4__bench;
	wire [0:0] n5_odata_p0_5__bench;
	wire [0:0] n5_odata_p0_6__bench;
	wire [0:0] n5_odata_p0_7__bench;
	wire [0:0] n5_odata_p0_8__bench;
	wire [0:0] n5_odata_p0_9__bench;
	wire [0:0] n5_odata_p0_10__bench;
	wire [0:0] n5_odata_p0_11__bench;
	wire [0:0] n5_odata_p0_12__bench;
	wire [0:0] n5_odata_p0_13__bench;
	wire [0:0] n5_odata_p0_14__bench;
	wire [0:0] n5_odata_p0_15__bench;
	wire [0:0] n5_odata_p0_16__bench;
	wire [0:0] n5_odata_p0_17__bench;
	wire [0:0] n5_odata_p0_18__bench;
	wire [0:0] n5_odata_p0_19__bench;
	wire [0:0] n5_odata_p0_20__bench;
	wire [0:0] n5_odata_p0_21__bench;
	wire [0:0] n5_odata_p0_22__bench;
	wire [0:0] n5_odata_p0_23__bench;
	wire [0:0] n5_odata_p0_24__bench;
	wire [0:0] n5_odata_p0_25__bench;
	wire [0:0] n5_odata_p0_26__bench;
	wire [0:0] n5_odata_p0_27__bench;
	wire [0:0] n5_odata_p0_28__bench;
	wire [0:0] n5_odata_p0_29__bench;
	wire [0:0] n5_odata_p0_30__bench;
	wire [0:0] n5_odata_p0_31__bench;
	wire [0:0] n5_odata_p0_32__bench;
	wire [0:0] n5_odata_p0_33__bench;
	wire [0:0] n5_odata_p0_34__bench;
	wire [0:0] n5_ovalid_p0_bench;
	wire [0:0] n6_ordy_p0_0__bench;
	wire [0:0] n6_ordy_p0_1__bench;
	wire [0:0] n6_odata_p0_0__bench;
	wire [0:0] n6_odata_p0_1__bench;
	wire [0:0] n6_odata_p0_2__bench;
	wire [0:0] n6_odata_p0_3__bench;
	wire [0:0] n6_odata_p0_4__bench;
	wire [0:0] n6_odata_p0_5__bench;
	wire [0:0] n6_odata_p0_6__bench;
	wire [0:0] n6_odata_p0_7__bench;
	wire [0:0] n6_odata_p0_8__bench;
	wire [0:0] n6_odata_p0_9__bench;
	wire [0:0] n6_odata_p0_10__bench;
	wire [0:0] n6_odata_p0_11__bench;
	wire [0:0] n6_odata_p0_12__bench;
	wire [0:0] n6_odata_p0_13__bench;
	wire [0:0] n6_odata_p0_14__bench;
	wire [0:0] n6_odata_p0_15__bench;
	wire [0:0] n6_odata_p0_16__bench;
	wire [0:0] n6_odata_p0_17__bench;
	wire [0:0] n6_odata_p0_18__bench;
	wire [0:0] n6_odata_p0_19__bench;
	wire [0:0] n6_odata_p0_20__bench;
	wire [0:0] n6_odata_p0_21__bench;
	wire [0:0] n6_odata_p0_22__bench;
	wire [0:0] n6_odata_p0_23__bench;
	wire [0:0] n6_odata_p0_24__bench;
	wire [0:0] n6_odata_p0_25__bench;
	wire [0:0] n6_odata_p0_26__bench;
	wire [0:0] n6_odata_p0_27__bench;
	wire [0:0] n6_odata_p0_28__bench;
	wire [0:0] n6_odata_p0_29__bench;
	wire [0:0] n6_odata_p0_30__bench;
	wire [0:0] n6_odata_p0_31__bench;
	wire [0:0] n6_odata_p0_32__bench;
	wire [0:0] n6_odata_p0_33__bench;
	wire [0:0] n6_odata_p0_34__bench;
	wire [0:0] n6_ovalid_p0_bench;
	wire [0:0] n7_ordy_p0_0__bench;
	wire [0:0] n7_ordy_p0_1__bench;
	wire [0:0] n7_odata_p0_0__bench;
	wire [0:0] n7_odata_p0_1__bench;
	wire [0:0] n7_odata_p0_2__bench;
	wire [0:0] n7_odata_p0_3__bench;
	wire [0:0] n7_odata_p0_4__bench;
	wire [0:0] n7_odata_p0_5__bench;
	wire [0:0] n7_odata_p0_6__bench;
	wire [0:0] n7_odata_p0_7__bench;
	wire [0:0] n7_odata_p0_8__bench;
	wire [0:0] n7_odata_p0_9__bench;
	wire [0:0] n7_odata_p0_10__bench;
	wire [0:0] n7_odata_p0_11__bench;
	wire [0:0] n7_odata_p0_12__bench;
	wire [0:0] n7_odata_p0_13__bench;
	wire [0:0] n7_odata_p0_14__bench;
	wire [0:0] n7_odata_p0_15__bench;
	wire [0:0] n7_odata_p0_16__bench;
	wire [0:0] n7_odata_p0_17__bench;
	wire [0:0] n7_odata_p0_18__bench;
	wire [0:0] n7_odata_p0_19__bench;
	wire [0:0] n7_odata_p0_20__bench;
	wire [0:0] n7_odata_p0_21__bench;
	wire [0:0] n7_odata_p0_22__bench;
	wire [0:0] n7_odata_p0_23__bench;
	wire [0:0] n7_odata_p0_24__bench;
	wire [0:0] n7_odata_p0_25__bench;
	wire [0:0] n7_odata_p0_26__bench;
	wire [0:0] n7_odata_p0_27__bench;
	wire [0:0] n7_odata_p0_28__bench;
	wire [0:0] n7_odata_p0_29__bench;
	wire [0:0] n7_odata_p0_30__bench;
	wire [0:0] n7_odata_p0_31__bench;
	wire [0:0] n7_odata_p0_32__bench;
	wire [0:0] n7_odata_p0_33__bench;
	wire [0:0] n7_odata_p0_34__bench;
	wire [0:0] n7_ovalid_p0_bench;
	wire [0:0] n8_ordy_p0_0__bench;
	wire [0:0] n8_ordy_p0_1__bench;
	wire [0:0] n8_odata_p0_0__bench;
	wire [0:0] n8_odata_p0_1__bench;
	wire [0:0] n8_odata_p0_2__bench;
	wire [0:0] n8_odata_p0_3__bench;
	wire [0:0] n8_odata_p0_4__bench;
	wire [0:0] n8_odata_p0_5__bench;
	wire [0:0] n8_odata_p0_6__bench;
	wire [0:0] n8_odata_p0_7__bench;
	wire [0:0] n8_odata_p0_8__bench;
	wire [0:0] n8_odata_p0_9__bench;
	wire [0:0] n8_odata_p0_10__bench;
	wire [0:0] n8_odata_p0_11__bench;
	wire [0:0] n8_odata_p0_12__bench;
	wire [0:0] n8_odata_p0_13__bench;
	wire [0:0] n8_odata_p0_14__bench;
	wire [0:0] n8_odata_p0_15__bench;
	wire [0:0] n8_odata_p0_16__bench;
	wire [0:0] n8_odata_p0_17__bench;
	wire [0:0] n8_odata_p0_18__bench;
	wire [0:0] n8_odata_p0_19__bench;
	wire [0:0] n8_odata_p0_20__bench;
	wire [0:0] n8_odata_p0_21__bench;
	wire [0:0] n8_odata_p0_22__bench;
	wire [0:0] n8_odata_p0_23__bench;
	wire [0:0] n8_odata_p0_24__bench;
	wire [0:0] n8_odata_p0_25__bench;
	wire [0:0] n8_odata_p0_26__bench;
	wire [0:0] n8_odata_p0_27__bench;
	wire [0:0] n8_odata_p0_28__bench;
	wire [0:0] n8_odata_p0_29__bench;
	wire [0:0] n8_odata_p0_30__bench;
	wire [0:0] n8_odata_p0_31__bench;
	wire [0:0] n8_odata_p0_32__bench;
	wire [0:0] n8_odata_p0_33__bench;
	wire [0:0] n8_odata_p0_34__bench;
	wire [0:0] n8_ovalid_p0_bench;

// ----- Output vectors checking flags -------
	reg [0:0] n0_ordy_p0_0__flag;
	reg [0:0] n0_ordy_p0_1__flag;
	reg [0:0] n0_odata_p0_0__flag;
	reg [0:0] n0_odata_p0_1__flag;
	reg [0:0] n0_odata_p0_2__flag;
	reg [0:0] n0_odata_p0_3__flag;
	reg [0:0] n0_odata_p0_4__flag;
	reg [0:0] n0_odata_p0_5__flag;
	reg [0:0] n0_odata_p0_6__flag;
	reg [0:0] n0_odata_p0_7__flag;
	reg [0:0] n0_odata_p0_8__flag;
	reg [0:0] n0_odata_p0_9__flag;
	reg [0:0] n0_odata_p0_10__flag;
	reg [0:0] n0_odata_p0_11__flag;
	reg [0:0] n0_odata_p0_12__flag;
	reg [0:0] n0_odata_p0_13__flag;
	reg [0:0] n0_odata_p0_14__flag;
	reg [0:0] n0_odata_p0_15__flag;
	reg [0:0] n0_odata_p0_16__flag;
	reg [0:0] n0_odata_p0_17__flag;
	reg [0:0] n0_odata_p0_18__flag;
	reg [0:0] n0_odata_p0_19__flag;
	reg [0:0] n0_odata_p0_20__flag;
	reg [0:0] n0_odata_p0_21__flag;
	reg [0:0] n0_odata_p0_22__flag;
	reg [0:0] n0_odata_p0_23__flag;
	reg [0:0] n0_odata_p0_24__flag;
	reg [0:0] n0_odata_p0_25__flag;
	reg [0:0] n0_odata_p0_26__flag;
	reg [0:0] n0_odata_p0_27__flag;
	reg [0:0] n0_odata_p0_28__flag;
	reg [0:0] n0_odata_p0_29__flag;
	reg [0:0] n0_odata_p0_30__flag;
	reg [0:0] n0_odata_p0_31__flag;
	reg [0:0] n0_odata_p0_32__flag;
	reg [0:0] n0_odata_p0_33__flag;
	reg [0:0] n0_odata_p0_34__flag;
	reg [0:0] n0_ovalid_p0_flag;
	reg [0:0] n1_ordy_p0_0__flag;
	reg [0:0] n1_ordy_p0_1__flag;
	reg [0:0] n1_odata_p0_0__flag;
	reg [0:0] n1_odata_p0_1__flag;
	reg [0:0] n1_odata_p0_2__flag;
	reg [0:0] n1_odata_p0_3__flag;
	reg [0:0] n1_odata_p0_4__flag;
	reg [0:0] n1_odata_p0_5__flag;
	reg [0:0] n1_odata_p0_6__flag;
	reg [0:0] n1_odata_p0_7__flag;
	reg [0:0] n1_odata_p0_8__flag;
	reg [0:0] n1_odata_p0_9__flag;
	reg [0:0] n1_odata_p0_10__flag;
	reg [0:0] n1_odata_p0_11__flag;
	reg [0:0] n1_odata_p0_12__flag;
	reg [0:0] n1_odata_p0_13__flag;
	reg [0:0] n1_odata_p0_14__flag;
	reg [0:0] n1_odata_p0_15__flag;
	reg [0:0] n1_odata_p0_16__flag;
	reg [0:0] n1_odata_p0_17__flag;
	reg [0:0] n1_odata_p0_18__flag;
	reg [0:0] n1_odata_p0_19__flag;
	reg [0:0] n1_odata_p0_20__flag;
	reg [0:0] n1_odata_p0_21__flag;
	reg [0:0] n1_odata_p0_22__flag;
	reg [0:0] n1_odata_p0_23__flag;
	reg [0:0] n1_odata_p0_24__flag;
	reg [0:0] n1_odata_p0_25__flag;
	reg [0:0] n1_odata_p0_26__flag;
	reg [0:0] n1_odata_p0_27__flag;
	reg [0:0] n1_odata_p0_28__flag;
	reg [0:0] n1_odata_p0_29__flag;
	reg [0:0] n1_odata_p0_30__flag;
	reg [0:0] n1_odata_p0_31__flag;
	reg [0:0] n1_odata_p0_32__flag;
	reg [0:0] n1_odata_p0_33__flag;
	reg [0:0] n1_odata_p0_34__flag;
	reg [0:0] n1_ovalid_p0_flag;
	reg [0:0] n2_ordy_p0_0__flag;
	reg [0:0] n2_ordy_p0_1__flag;
	reg [0:0] n2_odata_p0_0__flag;
	reg [0:0] n2_odata_p0_1__flag;
	reg [0:0] n2_odata_p0_2__flag;
	reg [0:0] n2_odata_p0_3__flag;
	reg [0:0] n2_odata_p0_4__flag;
	reg [0:0] n2_odata_p0_5__flag;
	reg [0:0] n2_odata_p0_6__flag;
	reg [0:0] n2_odata_p0_7__flag;
	reg [0:0] n2_odata_p0_8__flag;
	reg [0:0] n2_odata_p0_9__flag;
	reg [0:0] n2_odata_p0_10__flag;
	reg [0:0] n2_odata_p0_11__flag;
	reg [0:0] n2_odata_p0_12__flag;
	reg [0:0] n2_odata_p0_13__flag;
	reg [0:0] n2_odata_p0_14__flag;
	reg [0:0] n2_odata_p0_15__flag;
	reg [0:0] n2_odata_p0_16__flag;
	reg [0:0] n2_odata_p0_17__flag;
	reg [0:0] n2_odata_p0_18__flag;
	reg [0:0] n2_odata_p0_19__flag;
	reg [0:0] n2_odata_p0_20__flag;
	reg [0:0] n2_odata_p0_21__flag;
	reg [0:0] n2_odata_p0_22__flag;
	reg [0:0] n2_odata_p0_23__flag;
	reg [0:0] n2_odata_p0_24__flag;
	reg [0:0] n2_odata_p0_25__flag;
	reg [0:0] n2_odata_p0_26__flag;
	reg [0:0] n2_odata_p0_27__flag;
	reg [0:0] n2_odata_p0_28__flag;
	reg [0:0] n2_odata_p0_29__flag;
	reg [0:0] n2_odata_p0_30__flag;
	reg [0:0] n2_odata_p0_31__flag;
	reg [0:0] n2_odata_p0_32__flag;
	reg [0:0] n2_odata_p0_33__flag;
	reg [0:0] n2_odata_p0_34__flag;
	reg [0:0] n2_ovalid_p0_flag;
	reg [0:0] n3_ordy_p0_0__flag;
	reg [0:0] n3_ordy_p0_1__flag;
	reg [0:0] n3_odata_p0_0__flag;
	reg [0:0] n3_odata_p0_1__flag;
	reg [0:0] n3_odata_p0_2__flag;
	reg [0:0] n3_odata_p0_3__flag;
	reg [0:0] n3_odata_p0_4__flag;
	reg [0:0] n3_odata_p0_5__flag;
	reg [0:0] n3_odata_p0_6__flag;
	reg [0:0] n3_odata_p0_7__flag;
	reg [0:0] n3_odata_p0_8__flag;
	reg [0:0] n3_odata_p0_9__flag;
	reg [0:0] n3_odata_p0_10__flag;
	reg [0:0] n3_odata_p0_11__flag;
	reg [0:0] n3_odata_p0_12__flag;
	reg [0:0] n3_odata_p0_13__flag;
	reg [0:0] n3_odata_p0_14__flag;
	reg [0:0] n3_odata_p0_15__flag;
	reg [0:0] n3_odata_p0_16__flag;
	reg [0:0] n3_odata_p0_17__flag;
	reg [0:0] n3_odata_p0_18__flag;
	reg [0:0] n3_odata_p0_19__flag;
	reg [0:0] n3_odata_p0_20__flag;
	reg [0:0] n3_odata_p0_21__flag;
	reg [0:0] n3_odata_p0_22__flag;
	reg [0:0] n3_odata_p0_23__flag;
	reg [0:0] n3_odata_p0_24__flag;
	reg [0:0] n3_odata_p0_25__flag;
	reg [0:0] n3_odata_p0_26__flag;
	reg [0:0] n3_odata_p0_27__flag;
	reg [0:0] n3_odata_p0_28__flag;
	reg [0:0] n3_odata_p0_29__flag;
	reg [0:0] n3_odata_p0_30__flag;
	reg [0:0] n3_odata_p0_31__flag;
	reg [0:0] n3_odata_p0_32__flag;
	reg [0:0] n3_odata_p0_33__flag;
	reg [0:0] n3_odata_p0_34__flag;
	reg [0:0] n3_ovalid_p0_flag;
	reg [0:0] n4_ordy_p0_0__flag;
	reg [0:0] n4_ordy_p0_1__flag;
	reg [0:0] n4_odata_p0_0__flag;
	reg [0:0] n4_odata_p0_1__flag;
	reg [0:0] n4_odata_p0_2__flag;
	reg [0:0] n4_odata_p0_3__flag;
	reg [0:0] n4_odata_p0_4__flag;
	reg [0:0] n4_odata_p0_5__flag;
	reg [0:0] n4_odata_p0_6__flag;
	reg [0:0] n4_odata_p0_7__flag;
	reg [0:0] n4_odata_p0_8__flag;
	reg [0:0] n4_odata_p0_9__flag;
	reg [0:0] n4_odata_p0_10__flag;
	reg [0:0] n4_odata_p0_11__flag;
	reg [0:0] n4_odata_p0_12__flag;
	reg [0:0] n4_odata_p0_13__flag;
	reg [0:0] n4_odata_p0_14__flag;
	reg [0:0] n4_odata_p0_15__flag;
	reg [0:0] n4_odata_p0_16__flag;
	reg [0:0] n4_odata_p0_17__flag;
	reg [0:0] n4_odata_p0_18__flag;
	reg [0:0] n4_odata_p0_19__flag;
	reg [0:0] n4_odata_p0_20__flag;
	reg [0:0] n4_odata_p0_21__flag;
	reg [0:0] n4_odata_p0_22__flag;
	reg [0:0] n4_odata_p0_23__flag;
	reg [0:0] n4_odata_p0_24__flag;
	reg [0:0] n4_odata_p0_25__flag;
	reg [0:0] n4_odata_p0_26__flag;
	reg [0:0] n4_odata_p0_27__flag;
	reg [0:0] n4_odata_p0_28__flag;
	reg [0:0] n4_odata_p0_29__flag;
	reg [0:0] n4_odata_p0_30__flag;
	reg [0:0] n4_odata_p0_31__flag;
	reg [0:0] n4_odata_p0_32__flag;
	reg [0:0] n4_odata_p0_33__flag;
	reg [0:0] n4_odata_p0_34__flag;
	reg [0:0] n4_ovalid_p0_flag;
	reg [0:0] n5_ordy_p0_0__flag;
	reg [0:0] n5_ordy_p0_1__flag;
	reg [0:0] n5_odata_p0_0__flag;
	reg [0:0] n5_odata_p0_1__flag;
	reg [0:0] n5_odata_p0_2__flag;
	reg [0:0] n5_odata_p0_3__flag;
	reg [0:0] n5_odata_p0_4__flag;
	reg [0:0] n5_odata_p0_5__flag;
	reg [0:0] n5_odata_p0_6__flag;
	reg [0:0] n5_odata_p0_7__flag;
	reg [0:0] n5_odata_p0_8__flag;
	reg [0:0] n5_odata_p0_9__flag;
	reg [0:0] n5_odata_p0_10__flag;
	reg [0:0] n5_odata_p0_11__flag;
	reg [0:0] n5_odata_p0_12__flag;
	reg [0:0] n5_odata_p0_13__flag;
	reg [0:0] n5_odata_p0_14__flag;
	reg [0:0] n5_odata_p0_15__flag;
	reg [0:0] n5_odata_p0_16__flag;
	reg [0:0] n5_odata_p0_17__flag;
	reg [0:0] n5_odata_p0_18__flag;
	reg [0:0] n5_odata_p0_19__flag;
	reg [0:0] n5_odata_p0_20__flag;
	reg [0:0] n5_odata_p0_21__flag;
	reg [0:0] n5_odata_p0_22__flag;
	reg [0:0] n5_odata_p0_23__flag;
	reg [0:0] n5_odata_p0_24__flag;
	reg [0:0] n5_odata_p0_25__flag;
	reg [0:0] n5_odata_p0_26__flag;
	reg [0:0] n5_odata_p0_27__flag;
	reg [0:0] n5_odata_p0_28__flag;
	reg [0:0] n5_odata_p0_29__flag;
	reg [0:0] n5_odata_p0_30__flag;
	reg [0:0] n5_odata_p0_31__flag;
	reg [0:0] n5_odata_p0_32__flag;
	reg [0:0] n5_odata_p0_33__flag;
	reg [0:0] n5_odata_p0_34__flag;
	reg [0:0] n5_ovalid_p0_flag;
	reg [0:0] n6_ordy_p0_0__flag;
	reg [0:0] n6_ordy_p0_1__flag;
	reg [0:0] n6_odata_p0_0__flag;
	reg [0:0] n6_odata_p0_1__flag;
	reg [0:0] n6_odata_p0_2__flag;
	reg [0:0] n6_odata_p0_3__flag;
	reg [0:0] n6_odata_p0_4__flag;
	reg [0:0] n6_odata_p0_5__flag;
	reg [0:0] n6_odata_p0_6__flag;
	reg [0:0] n6_odata_p0_7__flag;
	reg [0:0] n6_odata_p0_8__flag;
	reg [0:0] n6_odata_p0_9__flag;
	reg [0:0] n6_odata_p0_10__flag;
	reg [0:0] n6_odata_p0_11__flag;
	reg [0:0] n6_odata_p0_12__flag;
	reg [0:0] n6_odata_p0_13__flag;
	reg [0:0] n6_odata_p0_14__flag;
	reg [0:0] n6_odata_p0_15__flag;
	reg [0:0] n6_odata_p0_16__flag;
	reg [0:0] n6_odata_p0_17__flag;
	reg [0:0] n6_odata_p0_18__flag;
	reg [0:0] n6_odata_p0_19__flag;
	reg [0:0] n6_odata_p0_20__flag;
	reg [0:0] n6_odata_p0_21__flag;
	reg [0:0] n6_odata_p0_22__flag;
	reg [0:0] n6_odata_p0_23__flag;
	reg [0:0] n6_odata_p0_24__flag;
	reg [0:0] n6_odata_p0_25__flag;
	reg [0:0] n6_odata_p0_26__flag;
	reg [0:0] n6_odata_p0_27__flag;
	reg [0:0] n6_odata_p0_28__flag;
	reg [0:0] n6_odata_p0_29__flag;
	reg [0:0] n6_odata_p0_30__flag;
	reg [0:0] n6_odata_p0_31__flag;
	reg [0:0] n6_odata_p0_32__flag;
	reg [0:0] n6_odata_p0_33__flag;
	reg [0:0] n6_odata_p0_34__flag;
	reg [0:0] n6_ovalid_p0_flag;
	reg [0:0] n7_ordy_p0_0__flag;
	reg [0:0] n7_ordy_p0_1__flag;
	reg [0:0] n7_odata_p0_0__flag;
	reg [0:0] n7_odata_p0_1__flag;
	reg [0:0] n7_odata_p0_2__flag;
	reg [0:0] n7_odata_p0_3__flag;
	reg [0:0] n7_odata_p0_4__flag;
	reg [0:0] n7_odata_p0_5__flag;
	reg [0:0] n7_odata_p0_6__flag;
	reg [0:0] n7_odata_p0_7__flag;
	reg [0:0] n7_odata_p0_8__flag;
	reg [0:0] n7_odata_p0_9__flag;
	reg [0:0] n7_odata_p0_10__flag;
	reg [0:0] n7_odata_p0_11__flag;
	reg [0:0] n7_odata_p0_12__flag;
	reg [0:0] n7_odata_p0_13__flag;
	reg [0:0] n7_odata_p0_14__flag;
	reg [0:0] n7_odata_p0_15__flag;
	reg [0:0] n7_odata_p0_16__flag;
	reg [0:0] n7_odata_p0_17__flag;
	reg [0:0] n7_odata_p0_18__flag;
	reg [0:0] n7_odata_p0_19__flag;
	reg [0:0] n7_odata_p0_20__flag;
	reg [0:0] n7_odata_p0_21__flag;
	reg [0:0] n7_odata_p0_22__flag;
	reg [0:0] n7_odata_p0_23__flag;
	reg [0:0] n7_odata_p0_24__flag;
	reg [0:0] n7_odata_p0_25__flag;
	reg [0:0] n7_odata_p0_26__flag;
	reg [0:0] n7_odata_p0_27__flag;
	reg [0:0] n7_odata_p0_28__flag;
	reg [0:0] n7_odata_p0_29__flag;
	reg [0:0] n7_odata_p0_30__flag;
	reg [0:0] n7_odata_p0_31__flag;
	reg [0:0] n7_odata_p0_32__flag;
	reg [0:0] n7_odata_p0_33__flag;
	reg [0:0] n7_odata_p0_34__flag;
	reg [0:0] n7_ovalid_p0_flag;
	reg [0:0] n8_ordy_p0_0__flag;
	reg [0:0] n8_ordy_p0_1__flag;
	reg [0:0] n8_odata_p0_0__flag;
	reg [0:0] n8_odata_p0_1__flag;
	reg [0:0] n8_odata_p0_2__flag;
	reg [0:0] n8_odata_p0_3__flag;
	reg [0:0] n8_odata_p0_4__flag;
	reg [0:0] n8_odata_p0_5__flag;
	reg [0:0] n8_odata_p0_6__flag;
	reg [0:0] n8_odata_p0_7__flag;
	reg [0:0] n8_odata_p0_8__flag;
	reg [0:0] n8_odata_p0_9__flag;
	reg [0:0] n8_odata_p0_10__flag;
	reg [0:0] n8_odata_p0_11__flag;
	reg [0:0] n8_odata_p0_12__flag;
	reg [0:0] n8_odata_p0_13__flag;
	reg [0:0] n8_odata_p0_14__flag;
	reg [0:0] n8_odata_p0_15__flag;
	reg [0:0] n8_odata_p0_16__flag;
	reg [0:0] n8_odata_p0_17__flag;
	reg [0:0] n8_odata_p0_18__flag;
	reg [0:0] n8_odata_p0_19__flag;
	reg [0:0] n8_odata_p0_20__flag;
	reg [0:0] n8_odata_p0_21__flag;
	reg [0:0] n8_odata_p0_22__flag;
	reg [0:0] n8_odata_p0_23__flag;
	reg [0:0] n8_odata_p0_24__flag;
	reg [0:0] n8_odata_p0_25__flag;
	reg [0:0] n8_odata_p0_26__flag;
	reg [0:0] n8_odata_p0_27__flag;
	reg [0:0] n8_odata_p0_28__flag;
	reg [0:0] n8_odata_p0_29__flag;
	reg [0:0] n8_odata_p0_30__flag;
	reg [0:0] n8_odata_p0_31__flag;
	reg [0:0] n8_odata_p0_32__flag;
	reg [0:0] n8_odata_p0_33__flag;
	reg [0:0] n8_odata_p0_34__flag;
	reg [0:0] n8_ovalid_p0_flag;

// ----- Error counter -------
	integer nb_error= 0;

// ----- FPGA fabric instanciation -------
	noc_top_formal_verification FPGA_DUT(
		n0_idata_p0_0_,
		n0_idata_p0_1_,
		n0_idata_p0_2_,
		n0_idata_p0_3_,
		n0_idata_p0_4_,
		n0_idata_p0_5_,
		n0_idata_p0_6_,
		n0_idata_p0_7_,
		n0_idata_p0_8_,
		n0_idata_p0_9_,
		n0_idata_p0_10_,
		n0_idata_p0_11_,
		n0_idata_p0_12_,
		n0_idata_p0_13_,
		n0_idata_p0_14_,
		n0_idata_p0_15_,
		n0_idata_p0_16_,
		n0_idata_p0_17_,
		n0_idata_p0_18_,
		n0_idata_p0_19_,
		n0_idata_p0_20_,
		n0_idata_p0_21_,
		n0_idata_p0_22_,
		n0_idata_p0_23_,
		n0_idata_p0_24_,
		n0_idata_p0_25_,
		n0_idata_p0_26_,
		n0_idata_p0_27_,
		n0_idata_p0_28_,
		n0_idata_p0_29_,
		n0_idata_p0_30_,
		n0_idata_p0_31_,
		n0_idata_p0_32_,
		n0_idata_p0_33_,
		n0_idata_p0_34_,
		n0_ivalid_p0,
		n0_ivch_p0,
		n1_idata_p0_0_,
		n1_idata_p0_1_,
		n1_idata_p0_2_,
		n1_idata_p0_3_,
		n1_idata_p0_4_,
		n1_idata_p0_5_,
		n1_idata_p0_6_,
		n1_idata_p0_7_,
		n1_idata_p0_8_,
		n1_idata_p0_9_,
		n1_idata_p0_10_,
		n1_idata_p0_11_,
		n1_idata_p0_12_,
		n1_idata_p0_13_,
		n1_idata_p0_14_,
		n1_idata_p0_15_,
		n1_idata_p0_16_,
		n1_idata_p0_17_,
		n1_idata_p0_18_,
		n1_idata_p0_19_,
		n1_idata_p0_20_,
		n1_idata_p0_21_,
		n1_idata_p0_22_,
		n1_idata_p0_23_,
		n1_idata_p0_24_,
		n1_idata_p0_25_,
		n1_idata_p0_26_,
		n1_idata_p0_27_,
		n1_idata_p0_28_,
		n1_idata_p0_29_,
		n1_idata_p0_30_,
		n1_idata_p0_31_,
		n1_idata_p0_32_,
		n1_idata_p0_33_,
		n1_idata_p0_34_,
		n1_ivalid_p0,
		n1_ivch_p0,
		n2_idata_p0_0_,
		n2_idata_p0_1_,
		n2_idata_p0_2_,
		n2_idata_p0_3_,
		n2_idata_p0_4_,
		n2_idata_p0_5_,
		n2_idata_p0_6_,
		n2_idata_p0_7_,
		n2_idata_p0_8_,
		n2_idata_p0_9_,
		n2_idata_p0_10_,
		n2_idata_p0_11_,
		n2_idata_p0_12_,
		n2_idata_p0_13_,
		n2_idata_p0_14_,
		n2_idata_p0_15_,
		n2_idata_p0_16_,
		n2_idata_p0_17_,
		n2_idata_p0_18_,
		n2_idata_p0_19_,
		n2_idata_p0_20_,
		n2_idata_p0_21_,
		n2_idata_p0_22_,
		n2_idata_p0_23_,
		n2_idata_p0_24_,
		n2_idata_p0_25_,
		n2_idata_p0_26_,
		n2_idata_p0_27_,
		n2_idata_p0_28_,
		n2_idata_p0_29_,
		n2_idata_p0_30_,
		n2_idata_p0_31_,
		n2_idata_p0_32_,
		n2_idata_p0_33_,
		n2_idata_p0_34_,
		n2_ivalid_p0,
		n2_ivch_p0,
		n3_idata_p0_0_,
		n3_idata_p0_1_,
		n3_idata_p0_2_,
		n3_idata_p0_3_,
		n3_idata_p0_4_,
		n3_idata_p0_5_,
		n3_idata_p0_6_,
		n3_idata_p0_7_,
		n3_idata_p0_8_,
		n3_idata_p0_9_,
		n3_idata_p0_10_,
		n3_idata_p0_11_,
		n3_idata_p0_12_,
		n3_idata_p0_13_,
		n3_idata_p0_14_,
		n3_idata_p0_15_,
		n3_idata_p0_16_,
		n3_idata_p0_17_,
		n3_idata_p0_18_,
		n3_idata_p0_19_,
		n3_idata_p0_20_,
		n3_idata_p0_21_,
		n3_idata_p0_22_,
		n3_idata_p0_23_,
		n3_idata_p0_24_,
		n3_idata_p0_25_,
		n3_idata_p0_26_,
		n3_idata_p0_27_,
		n3_idata_p0_28_,
		n3_idata_p0_29_,
		n3_idata_p0_30_,
		n3_idata_p0_31_,
		n3_idata_p0_32_,
		n3_idata_p0_33_,
		n3_idata_p0_34_,
		n3_ivalid_p0,
		n3_ivch_p0,
		n4_idata_p0_0_,
		n4_idata_p0_1_,
		n4_idata_p0_2_,
		n4_idata_p0_3_,
		n4_idata_p0_4_,
		n4_idata_p0_5_,
		n4_idata_p0_6_,
		n4_idata_p0_7_,
		n4_idata_p0_8_,
		n4_idata_p0_9_,
		n4_idata_p0_10_,
		n4_idata_p0_11_,
		n4_idata_p0_12_,
		n4_idata_p0_13_,
		n4_idata_p0_14_,
		n4_idata_p0_15_,
		n4_idata_p0_16_,
		n4_idata_p0_17_,
		n4_idata_p0_18_,
		n4_idata_p0_19_,
		n4_idata_p0_20_,
		n4_idata_p0_21_,
		n4_idata_p0_22_,
		n4_idata_p0_23_,
		n4_idata_p0_24_,
		n4_idata_p0_25_,
		n4_idata_p0_26_,
		n4_idata_p0_27_,
		n4_idata_p0_28_,
		n4_idata_p0_29_,
		n4_idata_p0_30_,
		n4_idata_p0_31_,
		n4_idata_p0_32_,
		n4_idata_p0_33_,
		n4_idata_p0_34_,
		n4_ivalid_p0,
		n4_ivch_p0,
		n5_idata_p0_0_,
		n5_idata_p0_1_,
		n5_idata_p0_2_,
		n5_idata_p0_3_,
		n5_idata_p0_4_,
		n5_idata_p0_5_,
		n5_idata_p0_6_,
		n5_idata_p0_7_,
		n5_idata_p0_8_,
		n5_idata_p0_9_,
		n5_idata_p0_10_,
		n5_idata_p0_11_,
		n5_idata_p0_12_,
		n5_idata_p0_13_,
		n5_idata_p0_14_,
		n5_idata_p0_15_,
		n5_idata_p0_16_,
		n5_idata_p0_17_,
		n5_idata_p0_18_,
		n5_idata_p0_19_,
		n5_idata_p0_20_,
		n5_idata_p0_21_,
		n5_idata_p0_22_,
		n5_idata_p0_23_,
		n5_idata_p0_24_,
		n5_idata_p0_25_,
		n5_idata_p0_26_,
		n5_idata_p0_27_,
		n5_idata_p0_28_,
		n5_idata_p0_29_,
		n5_idata_p0_30_,
		n5_idata_p0_31_,
		n5_idata_p0_32_,
		n5_idata_p0_33_,
		n5_idata_p0_34_,
		n5_ivalid_p0,
		n5_ivch_p0,
		n6_idata_p0_0_,
		n6_idata_p0_1_,
		n6_idata_p0_2_,
		n6_idata_p0_3_,
		n6_idata_p0_4_,
		n6_idata_p0_5_,
		n6_idata_p0_6_,
		n6_idata_p0_7_,
		n6_idata_p0_8_,
		n6_idata_p0_9_,
		n6_idata_p0_10_,
		n6_idata_p0_11_,
		n6_idata_p0_12_,
		n6_idata_p0_13_,
		n6_idata_p0_14_,
		n6_idata_p0_15_,
		n6_idata_p0_16_,
		n6_idata_p0_17_,
		n6_idata_p0_18_,
		n6_idata_p0_19_,
		n6_idata_p0_20_,
		n6_idata_p0_21_,
		n6_idata_p0_22_,
		n6_idata_p0_23_,
		n6_idata_p0_24_,
		n6_idata_p0_25_,
		n6_idata_p0_26_,
		n6_idata_p0_27_,
		n6_idata_p0_28_,
		n6_idata_p0_29_,
		n6_idata_p0_30_,
		n6_idata_p0_31_,
		n6_idata_p0_32_,
		n6_idata_p0_33_,
		n6_idata_p0_34_,
		n6_ivalid_p0,
		n6_ivch_p0,
		n7_idata_p0_0_,
		n7_idata_p0_1_,
		n7_idata_p0_2_,
		n7_idata_p0_3_,
		n7_idata_p0_4_,
		n7_idata_p0_5_,
		n7_idata_p0_6_,
		n7_idata_p0_7_,
		n7_idata_p0_8_,
		n7_idata_p0_9_,
		n7_idata_p0_10_,
		n7_idata_p0_11_,
		n7_idata_p0_12_,
		n7_idata_p0_13_,
		n7_idata_p0_14_,
		n7_idata_p0_15_,
		n7_idata_p0_16_,
		n7_idata_p0_17_,
		n7_idata_p0_18_,
		n7_idata_p0_19_,
		n7_idata_p0_20_,
		n7_idata_p0_21_,
		n7_idata_p0_22_,
		n7_idata_p0_23_,
		n7_idata_p0_24_,
		n7_idata_p0_25_,
		n7_idata_p0_26_,
		n7_idata_p0_27_,
		n7_idata_p0_28_,
		n7_idata_p0_29_,
		n7_idata_p0_30_,
		n7_idata_p0_31_,
		n7_idata_p0_32_,
		n7_idata_p0_33_,
		n7_idata_p0_34_,
		n7_ivalid_p0,
		n7_ivch_p0,
		n8_idata_p0_0_,
		n8_idata_p0_1_,
		n8_idata_p0_2_,
		n8_idata_p0_3_,
		n8_idata_p0_4_,
		n8_idata_p0_5_,
		n8_idata_p0_6_,
		n8_idata_p0_7_,
		n8_idata_p0_8_,
		n8_idata_p0_9_,
		n8_idata_p0_10_,
		n8_idata_p0_11_,
		n8_idata_p0_12_,
		n8_idata_p0_13_,
		n8_idata_p0_14_,
		n8_idata_p0_15_,
		n8_idata_p0_16_,
		n8_idata_p0_17_,
		n8_idata_p0_18_,
		n8_idata_p0_19_,
		n8_idata_p0_20_,
		n8_idata_p0_21_,
		n8_idata_p0_22_,
		n8_idata_p0_23_,
		n8_idata_p0_24_,
		n8_idata_p0_25_,
		n8_idata_p0_26_,
		n8_idata_p0_27_,
		n8_idata_p0_28_,
		n8_idata_p0_29_,
		n8_idata_p0_30_,
		n8_idata_p0_31_,
		n8_idata_p0_32_,
		n8_idata_p0_33_,
		n8_idata_p0_34_,
		n8_ivalid_p0,
		n8_ivch_p0,
		clk,
		rst_,
		n0_ordy_p0_0__gfpga,
		n0_ordy_p0_1__gfpga,
		n0_odata_p0_0__gfpga,
		n0_odata_p0_1__gfpga,
		n0_odata_p0_2__gfpga,
		n0_odata_p0_3__gfpga,
		n0_odata_p0_4__gfpga,
		n0_odata_p0_5__gfpga,
		n0_odata_p0_6__gfpga,
		n0_odata_p0_7__gfpga,
		n0_odata_p0_8__gfpga,
		n0_odata_p0_9__gfpga,
		n0_odata_p0_10__gfpga,
		n0_odata_p0_11__gfpga,
		n0_odata_p0_12__gfpga,
		n0_odata_p0_13__gfpga,
		n0_odata_p0_14__gfpga,
		n0_odata_p0_15__gfpga,
		n0_odata_p0_16__gfpga,
		n0_odata_p0_17__gfpga,
		n0_odata_p0_18__gfpga,
		n0_odata_p0_19__gfpga,
		n0_odata_p0_20__gfpga,
		n0_odata_p0_21__gfpga,
		n0_odata_p0_22__gfpga,
		n0_odata_p0_23__gfpga,
		n0_odata_p0_24__gfpga,
		n0_odata_p0_25__gfpga,
		n0_odata_p0_26__gfpga,
		n0_odata_p0_27__gfpga,
		n0_odata_p0_28__gfpga,
		n0_odata_p0_29__gfpga,
		n0_odata_p0_30__gfpga,
		n0_odata_p0_31__gfpga,
		n0_odata_p0_32__gfpga,
		n0_odata_p0_33__gfpga,
		n0_odata_p0_34__gfpga,
		n0_ovalid_p0_gfpga,
		n1_ordy_p0_0__gfpga,
		n1_ordy_p0_1__gfpga,
		n1_odata_p0_0__gfpga,
		n1_odata_p0_1__gfpga,
		n1_odata_p0_2__gfpga,
		n1_odata_p0_3__gfpga,
		n1_odata_p0_4__gfpga,
		n1_odata_p0_5__gfpga,
		n1_odata_p0_6__gfpga,
		n1_odata_p0_7__gfpga,
		n1_odata_p0_8__gfpga,
		n1_odata_p0_9__gfpga,
		n1_odata_p0_10__gfpga,
		n1_odata_p0_11__gfpga,
		n1_odata_p0_12__gfpga,
		n1_odata_p0_13__gfpga,
		n1_odata_p0_14__gfpga,
		n1_odata_p0_15__gfpga,
		n1_odata_p0_16__gfpga,
		n1_odata_p0_17__gfpga,
		n1_odata_p0_18__gfpga,
		n1_odata_p0_19__gfpga,
		n1_odata_p0_20__gfpga,
		n1_odata_p0_21__gfpga,
		n1_odata_p0_22__gfpga,
		n1_odata_p0_23__gfpga,
		n1_odata_p0_24__gfpga,
		n1_odata_p0_25__gfpga,
		n1_odata_p0_26__gfpga,
		n1_odata_p0_27__gfpga,
		n1_odata_p0_28__gfpga,
		n1_odata_p0_29__gfpga,
		n1_odata_p0_30__gfpga,
		n1_odata_p0_31__gfpga,
		n1_odata_p0_32__gfpga,
		n1_odata_p0_33__gfpga,
		n1_odata_p0_34__gfpga,
		n1_ovalid_p0_gfpga,
		n2_ordy_p0_0__gfpga,
		n2_ordy_p0_1__gfpga,
		n2_odata_p0_0__gfpga,
		n2_odata_p0_1__gfpga,
		n2_odata_p0_2__gfpga,
		n2_odata_p0_3__gfpga,
		n2_odata_p0_4__gfpga,
		n2_odata_p0_5__gfpga,
		n2_odata_p0_6__gfpga,
		n2_odata_p0_7__gfpga,
		n2_odata_p0_8__gfpga,
		n2_odata_p0_9__gfpga,
		n2_odata_p0_10__gfpga,
		n2_odata_p0_11__gfpga,
		n2_odata_p0_12__gfpga,
		n2_odata_p0_13__gfpga,
		n2_odata_p0_14__gfpga,
		n2_odata_p0_15__gfpga,
		n2_odata_p0_16__gfpga,
		n2_odata_p0_17__gfpga,
		n2_odata_p0_18__gfpga,
		n2_odata_p0_19__gfpga,
		n2_odata_p0_20__gfpga,
		n2_odata_p0_21__gfpga,
		n2_odata_p0_22__gfpga,
		n2_odata_p0_23__gfpga,
		n2_odata_p0_24__gfpga,
		n2_odata_p0_25__gfpga,
		n2_odata_p0_26__gfpga,
		n2_odata_p0_27__gfpga,
		n2_odata_p0_28__gfpga,
		n2_odata_p0_29__gfpga,
		n2_odata_p0_30__gfpga,
		n2_odata_p0_31__gfpga,
		n2_odata_p0_32__gfpga,
		n2_odata_p0_33__gfpga,
		n2_odata_p0_34__gfpga,
		n2_ovalid_p0_gfpga,
		n3_ordy_p0_0__gfpga,
		n3_ordy_p0_1__gfpga,
		n3_odata_p0_0__gfpga,
		n3_odata_p0_1__gfpga,
		n3_odata_p0_2__gfpga,
		n3_odata_p0_3__gfpga,
		n3_odata_p0_4__gfpga,
		n3_odata_p0_5__gfpga,
		n3_odata_p0_6__gfpga,
		n3_odata_p0_7__gfpga,
		n3_odata_p0_8__gfpga,
		n3_odata_p0_9__gfpga,
		n3_odata_p0_10__gfpga,
		n3_odata_p0_11__gfpga,
		n3_odata_p0_12__gfpga,
		n3_odata_p0_13__gfpga,
		n3_odata_p0_14__gfpga,
		n3_odata_p0_15__gfpga,
		n3_odata_p0_16__gfpga,
		n3_odata_p0_17__gfpga,
		n3_odata_p0_18__gfpga,
		n3_odata_p0_19__gfpga,
		n3_odata_p0_20__gfpga,
		n3_odata_p0_21__gfpga,
		n3_odata_p0_22__gfpga,
		n3_odata_p0_23__gfpga,
		n3_odata_p0_24__gfpga,
		n3_odata_p0_25__gfpga,
		n3_odata_p0_26__gfpga,
		n3_odata_p0_27__gfpga,
		n3_odata_p0_28__gfpga,
		n3_odata_p0_29__gfpga,
		n3_odata_p0_30__gfpga,
		n3_odata_p0_31__gfpga,
		n3_odata_p0_32__gfpga,
		n3_odata_p0_33__gfpga,
		n3_odata_p0_34__gfpga,
		n3_ovalid_p0_gfpga,
		n4_ordy_p0_0__gfpga,
		n4_ordy_p0_1__gfpga,
		n4_odata_p0_0__gfpga,
		n4_odata_p0_1__gfpga,
		n4_odata_p0_2__gfpga,
		n4_odata_p0_3__gfpga,
		n4_odata_p0_4__gfpga,
		n4_odata_p0_5__gfpga,
		n4_odata_p0_6__gfpga,
		n4_odata_p0_7__gfpga,
		n4_odata_p0_8__gfpga,
		n4_odata_p0_9__gfpga,
		n4_odata_p0_10__gfpga,
		n4_odata_p0_11__gfpga,
		n4_odata_p0_12__gfpga,
		n4_odata_p0_13__gfpga,
		n4_odata_p0_14__gfpga,
		n4_odata_p0_15__gfpga,
		n4_odata_p0_16__gfpga,
		n4_odata_p0_17__gfpga,
		n4_odata_p0_18__gfpga,
		n4_odata_p0_19__gfpga,
		n4_odata_p0_20__gfpga,
		n4_odata_p0_21__gfpga,
		n4_odata_p0_22__gfpga,
		n4_odata_p0_23__gfpga,
		n4_odata_p0_24__gfpga,
		n4_odata_p0_25__gfpga,
		n4_odata_p0_26__gfpga,
		n4_odata_p0_27__gfpga,
		n4_odata_p0_28__gfpga,
		n4_odata_p0_29__gfpga,
		n4_odata_p0_30__gfpga,
		n4_odata_p0_31__gfpga,
		n4_odata_p0_32__gfpga,
		n4_odata_p0_33__gfpga,
		n4_odata_p0_34__gfpga,
		n4_ovalid_p0_gfpga,
		n5_ordy_p0_0__gfpga,
		n5_ordy_p0_1__gfpga,
		n5_odata_p0_0__gfpga,
		n5_odata_p0_1__gfpga,
		n5_odata_p0_2__gfpga,
		n5_odata_p0_3__gfpga,
		n5_odata_p0_4__gfpga,
		n5_odata_p0_5__gfpga,
		n5_odata_p0_6__gfpga,
		n5_odata_p0_7__gfpga,
		n5_odata_p0_8__gfpga,
		n5_odata_p0_9__gfpga,
		n5_odata_p0_10__gfpga,
		n5_odata_p0_11__gfpga,
		n5_odata_p0_12__gfpga,
		n5_odata_p0_13__gfpga,
		n5_odata_p0_14__gfpga,
		n5_odata_p0_15__gfpga,
		n5_odata_p0_16__gfpga,
		n5_odata_p0_17__gfpga,
		n5_odata_p0_18__gfpga,
		n5_odata_p0_19__gfpga,
		n5_odata_p0_20__gfpga,
		n5_odata_p0_21__gfpga,
		n5_odata_p0_22__gfpga,
		n5_odata_p0_23__gfpga,
		n5_odata_p0_24__gfpga,
		n5_odata_p0_25__gfpga,
		n5_odata_p0_26__gfpga,
		n5_odata_p0_27__gfpga,
		n5_odata_p0_28__gfpga,
		n5_odata_p0_29__gfpga,
		n5_odata_p0_30__gfpga,
		n5_odata_p0_31__gfpga,
		n5_odata_p0_32__gfpga,
		n5_odata_p0_33__gfpga,
		n5_odata_p0_34__gfpga,
		n5_ovalid_p0_gfpga,
		n6_ordy_p0_0__gfpga,
		n6_ordy_p0_1__gfpga,
		n6_odata_p0_0__gfpga,
		n6_odata_p0_1__gfpga,
		n6_odata_p0_2__gfpga,
		n6_odata_p0_3__gfpga,
		n6_odata_p0_4__gfpga,
		n6_odata_p0_5__gfpga,
		n6_odata_p0_6__gfpga,
		n6_odata_p0_7__gfpga,
		n6_odata_p0_8__gfpga,
		n6_odata_p0_9__gfpga,
		n6_odata_p0_10__gfpga,
		n6_odata_p0_11__gfpga,
		n6_odata_p0_12__gfpga,
		n6_odata_p0_13__gfpga,
		n6_odata_p0_14__gfpga,
		n6_odata_p0_15__gfpga,
		n6_odata_p0_16__gfpga,
		n6_odata_p0_17__gfpga,
		n6_odata_p0_18__gfpga,
		n6_odata_p0_19__gfpga,
		n6_odata_p0_20__gfpga,
		n6_odata_p0_21__gfpga,
		n6_odata_p0_22__gfpga,
		n6_odata_p0_23__gfpga,
		n6_odata_p0_24__gfpga,
		n6_odata_p0_25__gfpga,
		n6_odata_p0_26__gfpga,
		n6_odata_p0_27__gfpga,
		n6_odata_p0_28__gfpga,
		n6_odata_p0_29__gfpga,
		n6_odata_p0_30__gfpga,
		n6_odata_p0_31__gfpga,
		n6_odata_p0_32__gfpga,
		n6_odata_p0_33__gfpga,
		n6_odata_p0_34__gfpga,
		n6_ovalid_p0_gfpga,
		n7_ordy_p0_0__gfpga,
		n7_ordy_p0_1__gfpga,
		n7_odata_p0_0__gfpga,
		n7_odata_p0_1__gfpga,
		n7_odata_p0_2__gfpga,
		n7_odata_p0_3__gfpga,
		n7_odata_p0_4__gfpga,
		n7_odata_p0_5__gfpga,
		n7_odata_p0_6__gfpga,
		n7_odata_p0_7__gfpga,
		n7_odata_p0_8__gfpga,
		n7_odata_p0_9__gfpga,
		n7_odata_p0_10__gfpga,
		n7_odata_p0_11__gfpga,
		n7_odata_p0_12__gfpga,
		n7_odata_p0_13__gfpga,
		n7_odata_p0_14__gfpga,
		n7_odata_p0_15__gfpga,
		n7_odata_p0_16__gfpga,
		n7_odata_p0_17__gfpga,
		n7_odata_p0_18__gfpga,
		n7_odata_p0_19__gfpga,
		n7_odata_p0_20__gfpga,
		n7_odata_p0_21__gfpga,
		n7_odata_p0_22__gfpga,
		n7_odata_p0_23__gfpga,
		n7_odata_p0_24__gfpga,
		n7_odata_p0_25__gfpga,
		n7_odata_p0_26__gfpga,
		n7_odata_p0_27__gfpga,
		n7_odata_p0_28__gfpga,
		n7_odata_p0_29__gfpga,
		n7_odata_p0_30__gfpga,
		n7_odata_p0_31__gfpga,
		n7_odata_p0_32__gfpga,
		n7_odata_p0_33__gfpga,
		n7_odata_p0_34__gfpga,
		n7_ovalid_p0_gfpga,
		n8_ordy_p0_0__gfpga,
		n8_ordy_p0_1__gfpga,
		n8_odata_p0_0__gfpga,
		n8_odata_p0_1__gfpga,
		n8_odata_p0_2__gfpga,
		n8_odata_p0_3__gfpga,
		n8_odata_p0_4__gfpga,
		n8_odata_p0_5__gfpga,
		n8_odata_p0_6__gfpga,
		n8_odata_p0_7__gfpga,
		n8_odata_p0_8__gfpga,
		n8_odata_p0_9__gfpga,
		n8_odata_p0_10__gfpga,
		n8_odata_p0_11__gfpga,
		n8_odata_p0_12__gfpga,
		n8_odata_p0_13__gfpga,
		n8_odata_p0_14__gfpga,
		n8_odata_p0_15__gfpga,
		n8_odata_p0_16__gfpga,
		n8_odata_p0_17__gfpga,
		n8_odata_p0_18__gfpga,
		n8_odata_p0_19__gfpga,
		n8_odata_p0_20__gfpga,
		n8_odata_p0_21__gfpga,
		n8_odata_p0_22__gfpga,
		n8_odata_p0_23__gfpga,
		n8_odata_p0_24__gfpga,
		n8_odata_p0_25__gfpga,
		n8_odata_p0_26__gfpga,
		n8_odata_p0_27__gfpga,
		n8_odata_p0_28__gfpga,
		n8_odata_p0_29__gfpga,
		n8_odata_p0_30__gfpga,
		n8_odata_p0_31__gfpga,
		n8_odata_p0_32__gfpga,
		n8_odata_p0_33__gfpga,
		n8_odata_p0_34__gfpga,
		n8_ovalid_p0_gfpga
	);
// ----- End FPGA Fabric Instanication -------

// ----- Reference Benchmark Instanication -------
	// noc REF_DUT(
	// 	n0_idata_p0_0_,
	// 	n0_idata_p0_1_,
	// 	n0_idata_p0_2_,
	// 	n0_idata_p0_3_,
	// 	n0_idata_p0_4_,
	// 	n0_idata_p0_5_,
	// 	n0_idata_p0_6_,
	// 	n0_idata_p0_7_,
	// 	n0_idata_p0_8_,
	// 	n0_idata_p0_9_,
	// 	n0_idata_p0_10_,
	// 	n0_idata_p0_11_,
	// 	n0_idata_p0_12_,
	// 	n0_idata_p0_13_,
	// 	n0_idata_p0_14_,
	// 	n0_idata_p0_15_,
	// 	n0_idata_p0_16_,
	// 	n0_idata_p0_17_,
	// 	n0_idata_p0_18_,
	// 	n0_idata_p0_19_,
	// 	n0_idata_p0_20_,
	// 	n0_idata_p0_21_,
	// 	n0_idata_p0_22_,
	// 	n0_idata_p0_23_,
	// 	n0_idata_p0_24_,
	// 	n0_idata_p0_25_,
	// 	n0_idata_p0_26_,
	// 	n0_idata_p0_27_,
	// 	n0_idata_p0_28_,
	// 	n0_idata_p0_29_,
	// 	n0_idata_p0_30_,
	// 	n0_idata_p0_31_,
	// 	n0_idata_p0_32_,
	// 	n0_idata_p0_33_,
	// 	n0_idata_p0_34_,
	// 	n0_ivalid_p0,
	// 	n0_ivch_p0,
	// 	n1_idata_p0_0_,
	// 	n1_idata_p0_1_,
	// 	n1_idata_p0_2_,
	// 	n1_idata_p0_3_,
	// 	n1_idata_p0_4_,
	// 	n1_idata_p0_5_,
	// 	n1_idata_p0_6_,
	// 	n1_idata_p0_7_,
	// 	n1_idata_p0_8_,
	// 	n1_idata_p0_9_,
	// 	n1_idata_p0_10_,
	// 	n1_idata_p0_11_,
	// 	n1_idata_p0_12_,
	// 	n1_idata_p0_13_,
	// 	n1_idata_p0_14_,
	// 	n1_idata_p0_15_,
	// 	n1_idata_p0_16_,
	// 	n1_idata_p0_17_,
	// 	n1_idata_p0_18_,
	// 	n1_idata_p0_19_,
	// 	n1_idata_p0_20_,
	// 	n1_idata_p0_21_,
	// 	n1_idata_p0_22_,
	// 	n1_idata_p0_23_,
	// 	n1_idata_p0_24_,
	// 	n1_idata_p0_25_,
	// 	n1_idata_p0_26_,
	// 	n1_idata_p0_27_,
	// 	n1_idata_p0_28_,
	// 	n1_idata_p0_29_,
	// 	n1_idata_p0_30_,
	// 	n1_idata_p0_31_,
	// 	n1_idata_p0_32_,
	// 	n1_idata_p0_33_,
	// 	n1_idata_p0_34_,
	// 	n1_ivalid_p0,
	// 	n1_ivch_p0,
	// 	n2_idata_p0_0_,
	// 	n2_idata_p0_1_,
	// 	n2_idata_p0_2_,
	// 	n2_idata_p0_3_,
	// 	n2_idata_p0_4_,
	// 	n2_idata_p0_5_,
	// 	n2_idata_p0_6_,
	// 	n2_idata_p0_7_,
	// 	n2_idata_p0_8_,
	// 	n2_idata_p0_9_,
	// 	n2_idata_p0_10_,
	// 	n2_idata_p0_11_,
	// 	n2_idata_p0_12_,
	// 	n2_idata_p0_13_,
	// 	n2_idata_p0_14_,
	// 	n2_idata_p0_15_,
	// 	n2_idata_p0_16_,
	// 	n2_idata_p0_17_,
	// 	n2_idata_p0_18_,
	// 	n2_idata_p0_19_,
	// 	n2_idata_p0_20_,
	// 	n2_idata_p0_21_,
	// 	n2_idata_p0_22_,
	// 	n2_idata_p0_23_,
	// 	n2_idata_p0_24_,
	// 	n2_idata_p0_25_,
	// 	n2_idata_p0_26_,
	// 	n2_idata_p0_27_,
	// 	n2_idata_p0_28_,
	// 	n2_idata_p0_29_,
	// 	n2_idata_p0_30_,
	// 	n2_idata_p0_31_,
	// 	n2_idata_p0_32_,
	// 	n2_idata_p0_33_,
	// 	n2_idata_p0_34_,
	// 	n2_ivalid_p0,
	// 	n2_ivch_p0,
	// 	n3_idata_p0_0_,
	// 	n3_idata_p0_1_,
	// 	n3_idata_p0_2_,
	// 	n3_idata_p0_3_,
	// 	n3_idata_p0_4_,
	// 	n3_idata_p0_5_,
	// 	n3_idata_p0_6_,
	// 	n3_idata_p0_7_,
	// 	n3_idata_p0_8_,
	// 	n3_idata_p0_9_,
	// 	n3_idata_p0_10_,
	// 	n3_idata_p0_11_,
	// 	n3_idata_p0_12_,
	// 	n3_idata_p0_13_,
	// 	n3_idata_p0_14_,
	// 	n3_idata_p0_15_,
	// 	n3_idata_p0_16_,
	// 	n3_idata_p0_17_,
	// 	n3_idata_p0_18_,
	// 	n3_idata_p0_19_,
	// 	n3_idata_p0_20_,
	// 	n3_idata_p0_21_,
	// 	n3_idata_p0_22_,
	// 	n3_idata_p0_23_,
	// 	n3_idata_p0_24_,
	// 	n3_idata_p0_25_,
	// 	n3_idata_p0_26_,
	// 	n3_idata_p0_27_,
	// 	n3_idata_p0_28_,
	// 	n3_idata_p0_29_,
	// 	n3_idata_p0_30_,
	// 	n3_idata_p0_31_,
	// 	n3_idata_p0_32_,
	// 	n3_idata_p0_33_,
	// 	n3_idata_p0_34_,
	// 	n3_ivalid_p0,
	// 	n3_ivch_p0,
	// 	n4_idata_p0_0_,
	// 	n4_idata_p0_1_,
	// 	n4_idata_p0_2_,
	// 	n4_idata_p0_3_,
	// 	n4_idata_p0_4_,
	// 	n4_idata_p0_5_,
	// 	n4_idata_p0_6_,
	// 	n4_idata_p0_7_,
	// 	n4_idata_p0_8_,
	// 	n4_idata_p0_9_,
	// 	n4_idata_p0_10_,
	// 	n4_idata_p0_11_,
	// 	n4_idata_p0_12_,
	// 	n4_idata_p0_13_,
	// 	n4_idata_p0_14_,
	// 	n4_idata_p0_15_,
	// 	n4_idata_p0_16_,
	// 	n4_idata_p0_17_,
	// 	n4_idata_p0_18_,
	// 	n4_idata_p0_19_,
	// 	n4_idata_p0_20_,
	// 	n4_idata_p0_21_,
	// 	n4_idata_p0_22_,
	// 	n4_idata_p0_23_,
	// 	n4_idata_p0_24_,
	// 	n4_idata_p0_25_,
	// 	n4_idata_p0_26_,
	// 	n4_idata_p0_27_,
	// 	n4_idata_p0_28_,
	// 	n4_idata_p0_29_,
	// 	n4_idata_p0_30_,
	// 	n4_idata_p0_31_,
	// 	n4_idata_p0_32_,
	// 	n4_idata_p0_33_,
	// 	n4_idata_p0_34_,
	// 	n4_ivalid_p0,
	// 	n4_ivch_p0,
	// 	n5_idata_p0_0_,
	// 	n5_idata_p0_1_,
	// 	n5_idata_p0_2_,
	// 	n5_idata_p0_3_,
	// 	n5_idata_p0_4_,
	// 	n5_idata_p0_5_,
	// 	n5_idata_p0_6_,
	// 	n5_idata_p0_7_,
	// 	n5_idata_p0_8_,
	// 	n5_idata_p0_9_,
	// 	n5_idata_p0_10_,
	// 	n5_idata_p0_11_,
	// 	n5_idata_p0_12_,
	// 	n5_idata_p0_13_,
	// 	n5_idata_p0_14_,
	// 	n5_idata_p0_15_,
	// 	n5_idata_p0_16_,
	// 	n5_idata_p0_17_,
	// 	n5_idata_p0_18_,
	// 	n5_idata_p0_19_,
	// 	n5_idata_p0_20_,
	// 	n5_idata_p0_21_,
	// 	n5_idata_p0_22_,
	// 	n5_idata_p0_23_,
	// 	n5_idata_p0_24_,
	// 	n5_idata_p0_25_,
	// 	n5_idata_p0_26_,
	// 	n5_idata_p0_27_,
	// 	n5_idata_p0_28_,
	// 	n5_idata_p0_29_,
	// 	n5_idata_p0_30_,
	// 	n5_idata_p0_31_,
	// 	n5_idata_p0_32_,
	// 	n5_idata_p0_33_,
	// 	n5_idata_p0_34_,
	// 	n5_ivalid_p0,
	// 	n5_ivch_p0,
	// 	n6_idata_p0_0_,
	// 	n6_idata_p0_1_,
	// 	n6_idata_p0_2_,
	// 	n6_idata_p0_3_,
	// 	n6_idata_p0_4_,
	// 	n6_idata_p0_5_,
	// 	n6_idata_p0_6_,
	// 	n6_idata_p0_7_,
	// 	n6_idata_p0_8_,
	// 	n6_idata_p0_9_,
	// 	n6_idata_p0_10_,
	// 	n6_idata_p0_11_,
	// 	n6_idata_p0_12_,
	// 	n6_idata_p0_13_,
	// 	n6_idata_p0_14_,
	// 	n6_idata_p0_15_,
	// 	n6_idata_p0_16_,
	// 	n6_idata_p0_17_,
	// 	n6_idata_p0_18_,
	// 	n6_idata_p0_19_,
	// 	n6_idata_p0_20_,
	// 	n6_idata_p0_21_,
	// 	n6_idata_p0_22_,
	// 	n6_idata_p0_23_,
	// 	n6_idata_p0_24_,
	// 	n6_idata_p0_25_,
	// 	n6_idata_p0_26_,
	// 	n6_idata_p0_27_,
	// 	n6_idata_p0_28_,
	// 	n6_idata_p0_29_,
	// 	n6_idata_p0_30_,
	// 	n6_idata_p0_31_,
	// 	n6_idata_p0_32_,
	// 	n6_idata_p0_33_,
	// 	n6_idata_p0_34_,
	// 	n6_ivalid_p0,
	// 	n6_ivch_p0,
	// 	n7_idata_p0_0_,
	// 	n7_idata_p0_1_,
	// 	n7_idata_p0_2_,
	// 	n7_idata_p0_3_,
	// 	n7_idata_p0_4_,
	// 	n7_idata_p0_5_,
	// 	n7_idata_p0_6_,
	// 	n7_idata_p0_7_,
	// 	n7_idata_p0_8_,
	// 	n7_idata_p0_9_,
	// 	n7_idata_p0_10_,
	// 	n7_idata_p0_11_,
	// 	n7_idata_p0_12_,
	// 	n7_idata_p0_13_,
	// 	n7_idata_p0_14_,
	// 	n7_idata_p0_15_,
	// 	n7_idata_p0_16_,
	// 	n7_idata_p0_17_,
	// 	n7_idata_p0_18_,
	// 	n7_idata_p0_19_,
	// 	n7_idata_p0_20_,
	// 	n7_idata_p0_21_,
	// 	n7_idata_p0_22_,
	// 	n7_idata_p0_23_,
	// 	n7_idata_p0_24_,
	// 	n7_idata_p0_25_,
	// 	n7_idata_p0_26_,
	// 	n7_idata_p0_27_,
	// 	n7_idata_p0_28_,
	// 	n7_idata_p0_29_,
	// 	n7_idata_p0_30_,
	// 	n7_idata_p0_31_,
	// 	n7_idata_p0_32_,
	// 	n7_idata_p0_33_,
	// 	n7_idata_p0_34_,
	// 	n7_ivalid_p0,
	// 	n7_ivch_p0,
	// 	n8_idata_p0_0_,
	// 	n8_idata_p0_1_,
	// 	n8_idata_p0_2_,
	// 	n8_idata_p0_3_,
	// 	n8_idata_p0_4_,
	// 	n8_idata_p0_5_,
	// 	n8_idata_p0_6_,
	// 	n8_idata_p0_7_,
	// 	n8_idata_p0_8_,
	// 	n8_idata_p0_9_,
	// 	n8_idata_p0_10_,
	// 	n8_idata_p0_11_,
	// 	n8_idata_p0_12_,
	// 	n8_idata_p0_13_,
	// 	n8_idata_p0_14_,
	// 	n8_idata_p0_15_,
	// 	n8_idata_p0_16_,
	// 	n8_idata_p0_17_,
	// 	n8_idata_p0_18_,
	// 	n8_idata_p0_19_,
	// 	n8_idata_p0_20_,
	// 	n8_idata_p0_21_,
	// 	n8_idata_p0_22_,
	// 	n8_idata_p0_23_,
	// 	n8_idata_p0_24_,
	// 	n8_idata_p0_25_,
	// 	n8_idata_p0_26_,
	// 	n8_idata_p0_27_,
	// 	n8_idata_p0_28_,
	// 	n8_idata_p0_29_,
	// 	n8_idata_p0_30_,
	// 	n8_idata_p0_31_,
	// 	n8_idata_p0_32_,
	// 	n8_idata_p0_33_,
	// 	n8_idata_p0_34_,
	// 	n8_ivalid_p0,
	// 	n8_ivch_p0,
	// 	clk,
	// 	rst_,
	// 	n0_ordy_p0_0__bench,
	// 	n0_ordy_p0_1__bench,
	// 	n0_odata_p0_0__bench,
	// 	n0_odata_p0_1__bench,
	// 	n0_odata_p0_2__bench,
	// 	n0_odata_p0_3__bench,
	// 	n0_odata_p0_4__bench,
	// 	n0_odata_p0_5__bench,
	// 	n0_odata_p0_6__bench,
	// 	n0_odata_p0_7__bench,
	// 	n0_odata_p0_8__bench,
	// 	n0_odata_p0_9__bench,
	// 	n0_odata_p0_10__bench,
	// 	n0_odata_p0_11__bench,
	// 	n0_odata_p0_12__bench,
	// 	n0_odata_p0_13__bench,
	// 	n0_odata_p0_14__bench,
	// 	n0_odata_p0_15__bench,
	// 	n0_odata_p0_16__bench,
	// 	n0_odata_p0_17__bench,
	// 	n0_odata_p0_18__bench,
	// 	n0_odata_p0_19__bench,
	// 	n0_odata_p0_20__bench,
	// 	n0_odata_p0_21__bench,
	// 	n0_odata_p0_22__bench,
	// 	n0_odata_p0_23__bench,
	// 	n0_odata_p0_24__bench,
	// 	n0_odata_p0_25__bench,
	// 	n0_odata_p0_26__bench,
	// 	n0_odata_p0_27__bench,
	// 	n0_odata_p0_28__bench,
	// 	n0_odata_p0_29__bench,
	// 	n0_odata_p0_30__bench,
	// 	n0_odata_p0_31__bench,
	// 	n0_odata_p0_32__bench,
	// 	n0_odata_p0_33__bench,
	// 	n0_odata_p0_34__bench,
	// 	n0_ovalid_p0_bench,
	// 	n1_ordy_p0_0__bench,
	// 	n1_ordy_p0_1__bench,
	// 	n1_odata_p0_0__bench,
	// 	n1_odata_p0_1__bench,
	// 	n1_odata_p0_2__bench,
	// 	n1_odata_p0_3__bench,
	// 	n1_odata_p0_4__bench,
	// 	n1_odata_p0_5__bench,
	// 	n1_odata_p0_6__bench,
	// 	n1_odata_p0_7__bench,
	// 	n1_odata_p0_8__bench,
	// 	n1_odata_p0_9__bench,
	// 	n1_odata_p0_10__bench,
	// 	n1_odata_p0_11__bench,
	// 	n1_odata_p0_12__bench,
	// 	n1_odata_p0_13__bench,
	// 	n1_odata_p0_14__bench,
	// 	n1_odata_p0_15__bench,
	// 	n1_odata_p0_16__bench,
	// 	n1_odata_p0_17__bench,
	// 	n1_odata_p0_18__bench,
	// 	n1_odata_p0_19__bench,
	// 	n1_odata_p0_20__bench,
	// 	n1_odata_p0_21__bench,
	// 	n1_odata_p0_22__bench,
	// 	n1_odata_p0_23__bench,
	// 	n1_odata_p0_24__bench,
	// 	n1_odata_p0_25__bench,
	// 	n1_odata_p0_26__bench,
	// 	n1_odata_p0_27__bench,
	// 	n1_odata_p0_28__bench,
	// 	n1_odata_p0_29__bench,
	// 	n1_odata_p0_30__bench,
	// 	n1_odata_p0_31__bench,
	// 	n1_odata_p0_32__bench,
	// 	n1_odata_p0_33__bench,
	// 	n1_odata_p0_34__bench,
	// 	n1_ovalid_p0_bench,
	// 	n2_ordy_p0_0__bench,
	// 	n2_ordy_p0_1__bench,
	// 	n2_odata_p0_0__bench,
	// 	n2_odata_p0_1__bench,
	// 	n2_odata_p0_2__bench,
	// 	n2_odata_p0_3__bench,
	// 	n2_odata_p0_4__bench,
	// 	n2_odata_p0_5__bench,
	// 	n2_odata_p0_6__bench,
	// 	n2_odata_p0_7__bench,
	// 	n2_odata_p0_8__bench,
	// 	n2_odata_p0_9__bench,
	// 	n2_odata_p0_10__bench,
	// 	n2_odata_p0_11__bench,
	// 	n2_odata_p0_12__bench,
	// 	n2_odata_p0_13__bench,
	// 	n2_odata_p0_14__bench,
	// 	n2_odata_p0_15__bench,
	// 	n2_odata_p0_16__bench,
	// 	n2_odata_p0_17__bench,
	// 	n2_odata_p0_18__bench,
	// 	n2_odata_p0_19__bench,
	// 	n2_odata_p0_20__bench,
	// 	n2_odata_p0_21__bench,
	// 	n2_odata_p0_22__bench,
	// 	n2_odata_p0_23__bench,
	// 	n2_odata_p0_24__bench,
	// 	n2_odata_p0_25__bench,
	// 	n2_odata_p0_26__bench,
	// 	n2_odata_p0_27__bench,
	// 	n2_odata_p0_28__bench,
	// 	n2_odata_p0_29__bench,
	// 	n2_odata_p0_30__bench,
	// 	n2_odata_p0_31__bench,
	// 	n2_odata_p0_32__bench,
	// 	n2_odata_p0_33__bench,
	// 	n2_odata_p0_34__bench,
	// 	n2_ovalid_p0_bench,
	// 	n3_ordy_p0_0__bench,
	// 	n3_ordy_p0_1__bench,
	// 	n3_odata_p0_0__bench,
	// 	n3_odata_p0_1__bench,
	// 	n3_odata_p0_2__bench,
	// 	n3_odata_p0_3__bench,
	// 	n3_odata_p0_4__bench,
	// 	n3_odata_p0_5__bench,
	// 	n3_odata_p0_6__bench,
	// 	n3_odata_p0_7__bench,
	// 	n3_odata_p0_8__bench,
	// 	n3_odata_p0_9__bench,
	// 	n3_odata_p0_10__bench,
	// 	n3_odata_p0_11__bench,
	// 	n3_odata_p0_12__bench,
	// 	n3_odata_p0_13__bench,
	// 	n3_odata_p0_14__bench,
	// 	n3_odata_p0_15__bench,
	// 	n3_odata_p0_16__bench,
	// 	n3_odata_p0_17__bench,
	// 	n3_odata_p0_18__bench,
	// 	n3_odata_p0_19__bench,
	// 	n3_odata_p0_20__bench,
	// 	n3_odata_p0_21__bench,
	// 	n3_odata_p0_22__bench,
	// 	n3_odata_p0_23__bench,
	// 	n3_odata_p0_24__bench,
	// 	n3_odata_p0_25__bench,
	// 	n3_odata_p0_26__bench,
	// 	n3_odata_p0_27__bench,
	// 	n3_odata_p0_28__bench,
	// 	n3_odata_p0_29__bench,
	// 	n3_odata_p0_30__bench,
	// 	n3_odata_p0_31__bench,
	// 	n3_odata_p0_32__bench,
	// 	n3_odata_p0_33__bench,
	// 	n3_odata_p0_34__bench,
	// 	n3_ovalid_p0_bench,
	// 	n4_ordy_p0_0__bench,
	// 	n4_ordy_p0_1__bench,
	// 	n4_odata_p0_0__bench,
	// 	n4_odata_p0_1__bench,
	// 	n4_odata_p0_2__bench,
	// 	n4_odata_p0_3__bench,
	// 	n4_odata_p0_4__bench,
	// 	n4_odata_p0_5__bench,
	// 	n4_odata_p0_6__bench,
	// 	n4_odata_p0_7__bench,
	// 	n4_odata_p0_8__bench,
	// 	n4_odata_p0_9__bench,
	// 	n4_odata_p0_10__bench,
	// 	n4_odata_p0_11__bench,
	// 	n4_odata_p0_12__bench,
	// 	n4_odata_p0_13__bench,
	// 	n4_odata_p0_14__bench,
	// 	n4_odata_p0_15__bench,
	// 	n4_odata_p0_16__bench,
	// 	n4_odata_p0_17__bench,
	// 	n4_odata_p0_18__bench,
	// 	n4_odata_p0_19__bench,
	// 	n4_odata_p0_20__bench,
	// 	n4_odata_p0_21__bench,
	// 	n4_odata_p0_22__bench,
	// 	n4_odata_p0_23__bench,
	// 	n4_odata_p0_24__bench,
	// 	n4_odata_p0_25__bench,
	// 	n4_odata_p0_26__bench,
	// 	n4_odata_p0_27__bench,
	// 	n4_odata_p0_28__bench,
	// 	n4_odata_p0_29__bench,
	// 	n4_odata_p0_30__bench,
	// 	n4_odata_p0_31__bench,
	// 	n4_odata_p0_32__bench,
	// 	n4_odata_p0_33__bench,
	// 	n4_odata_p0_34__bench,
	// 	n4_ovalid_p0_bench,
	// 	n5_ordy_p0_0__bench,
	// 	n5_ordy_p0_1__bench,
	// 	n5_odata_p0_0__bench,
	// 	n5_odata_p0_1__bench,
	// 	n5_odata_p0_2__bench,
	// 	n5_odata_p0_3__bench,
	// 	n5_odata_p0_4__bench,
	// 	n5_odata_p0_5__bench,
	// 	n5_odata_p0_6__bench,
	// 	n5_odata_p0_7__bench,
	// 	n5_odata_p0_8__bench,
	// 	n5_odata_p0_9__bench,
	// 	n5_odata_p0_10__bench,
	// 	n5_odata_p0_11__bench,
	// 	n5_odata_p0_12__bench,
	// 	n5_odata_p0_13__bench,
	// 	n5_odata_p0_14__bench,
	// 	n5_odata_p0_15__bench,
	// 	n5_odata_p0_16__bench,
	// 	n5_odata_p0_17__bench,
	// 	n5_odata_p0_18__bench,
	// 	n5_odata_p0_19__bench,
	// 	n5_odata_p0_20__bench,
	// 	n5_odata_p0_21__bench,
	// 	n5_odata_p0_22__bench,
	// 	n5_odata_p0_23__bench,
	// 	n5_odata_p0_24__bench,
	// 	n5_odata_p0_25__bench,
	// 	n5_odata_p0_26__bench,
	// 	n5_odata_p0_27__bench,
	// 	n5_odata_p0_28__bench,
	// 	n5_odata_p0_29__bench,
	// 	n5_odata_p0_30__bench,
	// 	n5_odata_p0_31__bench,
	// 	n5_odata_p0_32__bench,
	// 	n5_odata_p0_33__bench,
	// 	n5_odata_p0_34__bench,
	// 	n5_ovalid_p0_bench,
	// 	n6_ordy_p0_0__bench,
	// 	n6_ordy_p0_1__bench,
	// 	n6_odata_p0_0__bench,
	// 	n6_odata_p0_1__bench,
	// 	n6_odata_p0_2__bench,
	// 	n6_odata_p0_3__bench,
	// 	n6_odata_p0_4__bench,
	// 	n6_odata_p0_5__bench,
	// 	n6_odata_p0_6__bench,
	// 	n6_odata_p0_7__bench,
	// 	n6_odata_p0_8__bench,
	// 	n6_odata_p0_9__bench,
	// 	n6_odata_p0_10__bench,
	// 	n6_odata_p0_11__bench,
	// 	n6_odata_p0_12__bench,
	// 	n6_odata_p0_13__bench,
	// 	n6_odata_p0_14__bench,
	// 	n6_odata_p0_15__bench,
	// 	n6_odata_p0_16__bench,
	// 	n6_odata_p0_17__bench,
	// 	n6_odata_p0_18__bench,
	// 	n6_odata_p0_19__bench,
	// 	n6_odata_p0_20__bench,
	// 	n6_odata_p0_21__bench,
	// 	n6_odata_p0_22__bench,
	// 	n6_odata_p0_23__bench,
	// 	n6_odata_p0_24__bench,
	// 	n6_odata_p0_25__bench,
	// 	n6_odata_p0_26__bench,
	// 	n6_odata_p0_27__bench,
	// 	n6_odata_p0_28__bench,
	// 	n6_odata_p0_29__bench,
	// 	n6_odata_p0_30__bench,
	// 	n6_odata_p0_31__bench,
	// 	n6_odata_p0_32__bench,
	// 	n6_odata_p0_33__bench,
	// 	n6_odata_p0_34__bench,
	// 	n6_ovalid_p0_bench,
	// 	n7_ordy_p0_0__bench,
	// 	n7_ordy_p0_1__bench,
	// 	n7_odata_p0_0__bench,
	// 	n7_odata_p0_1__bench,
	// 	n7_odata_p0_2__bench,
	// 	n7_odata_p0_3__bench,
	// 	n7_odata_p0_4__bench,
	// 	n7_odata_p0_5__bench,
	// 	n7_odata_p0_6__bench,
	// 	n7_odata_p0_7__bench,
	// 	n7_odata_p0_8__bench,
	// 	n7_odata_p0_9__bench,
	// 	n7_odata_p0_10__bench,
	// 	n7_odata_p0_11__bench,
	// 	n7_odata_p0_12__bench,
	// 	n7_odata_p0_13__bench,
	// 	n7_odata_p0_14__bench,
	// 	n7_odata_p0_15__bench,
	// 	n7_odata_p0_16__bench,
	// 	n7_odata_p0_17__bench,
	// 	n7_odata_p0_18__bench,
	// 	n7_odata_p0_19__bench,
	// 	n7_odata_p0_20__bench,
	// 	n7_odata_p0_21__bench,
	// 	n7_odata_p0_22__bench,
	// 	n7_odata_p0_23__bench,
	// 	n7_odata_p0_24__bench,
	// 	n7_odata_p0_25__bench,
	// 	n7_odata_p0_26__bench,
	// 	n7_odata_p0_27__bench,
	// 	n7_odata_p0_28__bench,
	// 	n7_odata_p0_29__bench,
	// 	n7_odata_p0_30__bench,
	// 	n7_odata_p0_31__bench,
	// 	n7_odata_p0_32__bench,
	// 	n7_odata_p0_33__bench,
	// 	n7_odata_p0_34__bench,
	// 	n7_ovalid_p0_bench,
	// 	n8_ordy_p0_0__bench,
	// 	n8_ordy_p0_1__bench,
	// 	n8_odata_p0_0__bench,
	// 	n8_odata_p0_1__bench,
	// 	n8_odata_p0_2__bench,
	// 	n8_odata_p0_3__bench,
	// 	n8_odata_p0_4__bench,
	// 	n8_odata_p0_5__bench,
	// 	n8_odata_p0_6__bench,
	// 	n8_odata_p0_7__bench,
	// 	n8_odata_p0_8__bench,
	// 	n8_odata_p0_9__bench,
	// 	n8_odata_p0_10__bench,
	// 	n8_odata_p0_11__bench,
	// 	n8_odata_p0_12__bench,
	// 	n8_odata_p0_13__bench,
	// 	n8_odata_p0_14__bench,
	// 	n8_odata_p0_15__bench,
	// 	n8_odata_p0_16__bench,
	// 	n8_odata_p0_17__bench,
	// 	n8_odata_p0_18__bench,
	// 	n8_odata_p0_19__bench,
	// 	n8_odata_p0_20__bench,
	// 	n8_odata_p0_21__bench,
	// 	n8_odata_p0_22__bench,
	// 	n8_odata_p0_23__bench,
	// 	n8_odata_p0_24__bench,
	// 	n8_odata_p0_25__bench,
	// 	n8_odata_p0_26__bench,
	// 	n8_odata_p0_27__bench,
	// 	n8_odata_p0_28__bench,
	// 	n8_odata_p0_29__bench,
	// 	n8_odata_p0_30__bench,
	// 	n8_odata_p0_31__bench,
	// 	n8_odata_p0_32__bench,
	// 	n8_odata_p0_33__bench,
	// 	n8_odata_p0_34__bench,
	// 	n8_ovalid_p0_bench
	// );

	noc REF_DUT(
		.n0_idata_p0({n0_idata_p0_0_,
		n0_idata_p0_1_,
		n0_idata_p0_2_,
		n0_idata_p0_3_,
		n0_idata_p0_4_,
		n0_idata_p0_5_,
		n0_idata_p0_6_,
		n0_idata_p0_7_,
		n0_idata_p0_8_,
		n0_idata_p0_9_,
		n0_idata_p0_10_,
		n0_idata_p0_11_,
		n0_idata_p0_12_,
		n0_idata_p0_13_,
		n0_idata_p0_14_,
		n0_idata_p0_15_,
		n0_idata_p0_16_,
		n0_idata_p0_17_,
		n0_idata_p0_18_,
		n0_idata_p0_19_,
		n0_idata_p0_20_,
		n0_idata_p0_21_,
		n0_idata_p0_22_,
		n0_idata_p0_23_,
		n0_idata_p0_24_,
		n0_idata_p0_25_,
		n0_idata_p0_26_,
		n0_idata_p0_27_,
		n0_idata_p0_28_,
		n0_idata_p0_29_,
		n0_idata_p0_30_,
		n0_idata_p0_31_,
		n0_idata_p0_32_,
		n0_idata_p0_33_,
		n0_idata_p0_34_}),
		.n0_ivalid_p0(n0_ivalid_p0),
		.n0_ivch_p0(n0_ivch_p0),
		.n1_idata_p0({n1_idata_p0_0_,
		n1_idata_p0_1_,
		n1_idata_p0_2_,
		n1_idata_p0_3_,
		n1_idata_p0_4_,
		n1_idata_p0_5_,
		n1_idata_p0_6_,
		n1_idata_p0_7_,
		n1_idata_p0_8_,
		n1_idata_p0_9_,
		n1_idata_p0_10_,
		n1_idata_p0_11_,
		n1_idata_p0_12_,
		n1_idata_p0_13_,
		n1_idata_p0_14_,
		n1_idata_p0_15_,
		n1_idata_p0_16_,
		n1_idata_p0_17_,
		n1_idata_p0_18_,
		n1_idata_p0_19_,
		n1_idata_p0_20_,
		n1_idata_p0_21_,
		n1_idata_p0_22_,
		n1_idata_p0_23_,
		n1_idata_p0_24_,
		n1_idata_p0_25_,
		n1_idata_p0_26_,
		n1_idata_p0_27_,
		n1_idata_p0_28_,
		n1_idata_p0_29_,
		n1_idata_p0_30_,
		n1_idata_p0_31_,
		n1_idata_p0_32_,
		n1_idata_p0_33_,
		n1_idata_p0_34_}),
		.n1_ivalid_p0(n1_ivalid_p0),
		.n1_ivch_p0(n1_ivch_p0),
		.n2_idata_p0({n2_idata_p0_0_,
		n2_idata_p0_1_,
		n2_idata_p0_2_,
		n2_idata_p0_3_,
		n2_idata_p0_4_,
		n2_idata_p0_5_,
		n2_idata_p0_6_,
		n2_idata_p0_7_,
		n2_idata_p0_8_,
		n2_idata_p0_9_,
		n2_idata_p0_10_,
		n2_idata_p0_11_,
		n2_idata_p0_12_,
		n2_idata_p0_13_,
		n2_idata_p0_14_,
		n2_idata_p0_15_,
		n2_idata_p0_16_,
		n2_idata_p0_17_,
		n2_idata_p0_18_,
		n2_idata_p0_19_,
		n2_idata_p0_20_,
		n2_idata_p0_21_,
		n2_idata_p0_22_,
		n2_idata_p0_23_,
		n2_idata_p0_24_,
		n2_idata_p0_25_,
		n2_idata_p0_26_,
		n2_idata_p0_27_,
		n2_idata_p0_28_,
		n2_idata_p0_29_,
		n2_idata_p0_30_,
		n2_idata_p0_31_,
		n2_idata_p0_32_,
		n2_idata_p0_33_,
		n2_idata_p0_34_}),
		.n2_ivalid_p0(n2_ivalid_p0),
		.n2_ivch_p0(n2_ivch_p0),
		.n3_idata_p0({n3_idata_p0_0_,
		n3_idata_p0_1_,
		n3_idata_p0_2_,
		n3_idata_p0_3_,
		n3_idata_p0_4_,
		n3_idata_p0_5_,
		n3_idata_p0_6_,
		n3_idata_p0_7_,
		n3_idata_p0_8_,
		n3_idata_p0_9_,
		n3_idata_p0_10_,
		n3_idata_p0_11_,
		n3_idata_p0_12_,
		n3_idata_p0_13_,
		n3_idata_p0_14_,
		n3_idata_p0_15_,
		n3_idata_p0_16_,
		n3_idata_p0_17_,
		n3_idata_p0_18_,
		n3_idata_p0_19_,
		n3_idata_p0_20_,
		n3_idata_p0_21_,
		n3_idata_p0_22_,
		n3_idata_p0_23_,
		n3_idata_p0_24_,
		n3_idata_p0_25_,
		n3_idata_p0_26_,
		n3_idata_p0_27_,
		n3_idata_p0_28_,
		n3_idata_p0_29_,
		n3_idata_p0_30_,
		n3_idata_p0_31_,
		n3_idata_p0_32_,
		n3_idata_p0_33_,
		n3_idata_p0_34_}),
		.n3_ivalid_p0(n3_ivalid_p0),
		.n3_ivch_p0(n3_ivch_p0),
		.n4_idata_p0({n4_idata_p0_0_,
		n4_idata_p0_1_,
		n4_idata_p0_2_,
		n4_idata_p0_3_,
		n4_idata_p0_4_,
		n4_idata_p0_5_,
		n4_idata_p0_6_,
		n4_idata_p0_7_,
		n4_idata_p0_8_,
		n4_idata_p0_9_,
		n4_idata_p0_10_,
		n4_idata_p0_11_,
		n4_idata_p0_12_,
		n4_idata_p0_13_,
		n4_idata_p0_14_,
		n4_idata_p0_15_,
		n4_idata_p0_16_,
		n4_idata_p0_17_,
		n4_idata_p0_18_,
		n4_idata_p0_19_,
		n4_idata_p0_20_,
		n4_idata_p0_21_,
		n4_idata_p0_22_,
		n4_idata_p0_23_,
		n4_idata_p0_24_,
		n4_idata_p0_25_,
		n4_idata_p0_26_,
		n4_idata_p0_27_,
		n4_idata_p0_28_,
		n4_idata_p0_29_,
		n4_idata_p0_30_,
		n4_idata_p0_31_,
		n4_idata_p0_32_,
		n4_idata_p0_33_,
		n4_idata_p0_34_}),
		.n4_ivalid_p0(n4_ivalid_p0),
		.n4_ivch_p0(n4_ivch_p0),
		.n5_idata_p0({n5_idata_p0_0_,
		n5_idata_p0_1_,
		n5_idata_p0_2_,
		n5_idata_p0_3_,
		n5_idata_p0_4_,
		n5_idata_p0_5_,
		n5_idata_p0_6_,
		n5_idata_p0_7_,
		n5_idata_p0_8_,
		n5_idata_p0_9_,
		n5_idata_p0_10_,
		n5_idata_p0_11_,
		n5_idata_p0_12_,
		n5_idata_p0_13_,
		n5_idata_p0_14_,
		n5_idata_p0_15_,
		n5_idata_p0_16_,
		n5_idata_p0_17_,
		n5_idata_p0_18_,
		n5_idata_p0_19_,
		n5_idata_p0_20_,
		n5_idata_p0_21_,
		n5_idata_p0_22_,
		n5_idata_p0_23_,
		n5_idata_p0_24_,
		n5_idata_p0_25_,
		n5_idata_p0_26_,
		n5_idata_p0_27_,
		n5_idata_p0_28_,
		n5_idata_p0_29_,
		n5_idata_p0_30_,
		n5_idata_p0_31_,
		n5_idata_p0_32_,
		n5_idata_p0_33_,
		n5_idata_p0_34_}),
		.n5_ivalid_p0(n5_ivalid_p0),
		.n5_ivch_p0(n5_ivch_p0),
		.n6_idata_p0({n6_idata_p0_0_,
		n6_idata_p0_1_,
		n6_idata_p0_2_,
		n6_idata_p0_3_,
		n6_idata_p0_4_,
		n6_idata_p0_5_,
		n6_idata_p0_6_,
		n6_idata_p0_7_,
		n6_idata_p0_8_,
		n6_idata_p0_9_,
		n6_idata_p0_10_,
		n6_idata_p0_11_,
		n6_idata_p0_12_,
		n6_idata_p0_13_,
		n6_idata_p0_14_,
		n6_idata_p0_15_,
		n6_idata_p0_16_,
		n6_idata_p0_17_,
		n6_idata_p0_18_,
		n6_idata_p0_19_,
		n6_idata_p0_20_,
		n6_idata_p0_21_,
		n6_idata_p0_22_,
		n6_idata_p0_23_,
		n6_idata_p0_24_,
		n6_idata_p0_25_,
		n6_idata_p0_26_,
		n6_idata_p0_27_,
		n6_idata_p0_28_,
		n6_idata_p0_29_,
		n6_idata_p0_30_,
		n6_idata_p0_31_,
		n6_idata_p0_32_,
		n6_idata_p0_33_,
		n6_idata_p0_34_}),
		.n6_ivalid_p0(n6_ivalid_p0),
		.n6_ivch_p0(n6_ivch_p0),
		.n7_idata_p0({n7_idata_p0_0_,
		n7_idata_p0_1_,
		n7_idata_p0_2_,
		n7_idata_p0_3_,
		n7_idata_p0_4_,
		n7_idata_p0_5_,
		n7_idata_p0_6_,
		n7_idata_p0_7_,
		n7_idata_p0_8_,
		n7_idata_p0_9_,
		n7_idata_p0_10_,
		n7_idata_p0_11_,
		n7_idata_p0_12_,
		n7_idata_p0_13_,
		n7_idata_p0_14_,
		n7_idata_p0_15_,
		n7_idata_p0_16_,
		n7_idata_p0_17_,
		n7_idata_p0_18_,
		n7_idata_p0_19_,
		n7_idata_p0_20_,
		n7_idata_p0_21_,
		n7_idata_p0_22_,
		n7_idata_p0_23_,
		n7_idata_p0_24_,
		n7_idata_p0_25_,
		n7_idata_p0_26_,
		n7_idata_p0_27_,
		n7_idata_p0_28_,
		n7_idata_p0_29_,
		n7_idata_p0_30_,
		n7_idata_p0_31_,
		n7_idata_p0_32_,
		n7_idata_p0_33_,
		n7_idata_p0_34_}),
		.n7_ivalid_p0(n7_ivalid_p0),
		.n7_ivch_p0(n7_ivch_p0),
		.n8_idata_p0({n8_idata_p0_0_,
		n8_idata_p0_1_,
		n8_idata_p0_2_,
		n8_idata_p0_3_,
		n8_idata_p0_4_,
		n8_idata_p0_5_,
		n8_idata_p0_6_,
		n8_idata_p0_7_,
		n8_idata_p0_8_,
		n8_idata_p0_9_,
		n8_idata_p0_10_,
		n8_idata_p0_11_,
		n8_idata_p0_12_,
		n8_idata_p0_13_,
		n8_idata_p0_14_,
		n8_idata_p0_15_,
		n8_idata_p0_16_,
		n8_idata_p0_17_,
		n8_idata_p0_18_,
		n8_idata_p0_19_,
		n8_idata_p0_20_,
		n8_idata_p0_21_,
		n8_idata_p0_22_,
		n8_idata_p0_23_,
		n8_idata_p0_24_,
		n8_idata_p0_25_,
		n8_idata_p0_26_,
		n8_idata_p0_27_,
		n8_idata_p0_28_,
		n8_idata_p0_29_,
		n8_idata_p0_30_,
		n8_idata_p0_31_,
		n8_idata_p0_32_,
		n8_idata_p0_33_,
		n8_idata_p0_34_}),
		.n8_ivalid_p0(n8_ivalid_p0),
		.n8_ivch_p0(n8_ivch_p0),
		.clk(clk),
		.rst_(rst_),
		.n0_ordy_p0({n0_ordy_p0_0__bench,
		n0_ordy_p0_1__bench}),
		.n0_odata_p0({n0_odata_p0_0__bench,
		n0_odata_p0_1__bench,
		n0_odata_p0_2__bench,
		n0_odata_p0_3__bench,
		n0_odata_p0_4__bench,
		n0_odata_p0_5__bench,
		n0_odata_p0_6__bench,
		n0_odata_p0_7__bench,
		n0_odata_p0_8__bench,
		n0_odata_p0_9__bench,
		n0_odata_p0_10__bench,
		n0_odata_p0_11__bench,
		n0_odata_p0_12__bench,
		n0_odata_p0_13__bench,
		n0_odata_p0_14__bench,
		n0_odata_p0_15__bench,
		n0_odata_p0_16__bench,
		n0_odata_p0_17__bench,
		n0_odata_p0_18__bench,
		n0_odata_p0_19__bench,
		n0_odata_p0_20__bench,
		n0_odata_p0_21__bench,
		n0_odata_p0_22__bench,
		n0_odata_p0_23__bench,
		n0_odata_p0_24__bench,
		n0_odata_p0_25__bench,
		n0_odata_p0_26__bench,
		n0_odata_p0_27__bench,
		n0_odata_p0_28__bench,
		n0_odata_p0_29__bench,
		n0_odata_p0_30__bench,
		n0_odata_p0_31__bench,
		n0_odata_p0_32__bench,
		n0_odata_p0_33__bench,
		n0_odata_p0_34__bench}),
		.n0_ovalid_p0({n0_ovalid_p0_bench}),
		.n1_ordy_p0({n1_ordy_p0_0__bench,
		n1_ordy_p0_1__bench}),
		.n1_odata_p0({n1_odata_p0_0__bench,
		n1_odata_p0_1__bench,
		n1_odata_p0_2__bench,
		n1_odata_p0_3__bench,
		n1_odata_p0_4__bench,
		n1_odata_p0_5__bench,
		n1_odata_p0_6__bench,
		n1_odata_p0_7__bench,
		n1_odata_p0_8__bench,
		n1_odata_p0_9__bench,
		n1_odata_p0_10__bench,
		n1_odata_p0_11__bench,
		n1_odata_p0_12__bench,
		n1_odata_p0_13__bench,
		n1_odata_p0_14__bench,
		n1_odata_p0_15__bench,
		n1_odata_p0_16__bench,
		n1_odata_p0_17__bench,
		n1_odata_p0_18__bench,
		n1_odata_p0_19__bench,
		n1_odata_p0_20__bench,
		n1_odata_p0_21__bench,
		n1_odata_p0_22__bench,
		n1_odata_p0_23__bench,
		n1_odata_p0_24__bench,
		n1_odata_p0_25__bench,
		n1_odata_p0_26__bench,
		n1_odata_p0_27__bench,
		n1_odata_p0_28__bench,
		n1_odata_p0_29__bench,
		n1_odata_p0_30__bench,
		n1_odata_p0_31__bench,
		n1_odata_p0_32__bench,
		n1_odata_p0_33__bench,
		n1_odata_p0_34__bench}),
		.n1_ovalid_p0(n1_ovalid_p0_bench),
		.n2_ordy_p0({n2_ordy_p0_0__bench,
		n2_ordy_p0_1__bench}),
		.n2_odata_p0({n2_odata_p0_0__bench,
		n2_odata_p0_1__bench,
		n2_odata_p0_2__bench,
		n2_odata_p0_3__bench,
		n2_odata_p0_4__bench,
		n2_odata_p0_5__bench,
		n2_odata_p0_6__bench,
		n2_odata_p0_7__bench,
		n2_odata_p0_8__bench,
		n2_odata_p0_9__bench,
		n2_odata_p0_10__bench,
		n2_odata_p0_11__bench,
		n2_odata_p0_12__bench,
		n2_odata_p0_13__bench,
		n2_odata_p0_14__bench,
		n2_odata_p0_15__bench,
		n2_odata_p0_16__bench,
		n2_odata_p0_17__bench,
		n2_odata_p0_18__bench,
		n2_odata_p0_19__bench,
		n2_odata_p0_20__bench,
		n2_odata_p0_21__bench,
		n2_odata_p0_22__bench,
		n2_odata_p0_23__bench,
		n2_odata_p0_24__bench,
		n2_odata_p0_25__bench,
		n2_odata_p0_26__bench,
		n2_odata_p0_27__bench,
		n2_odata_p0_28__bench,
		n2_odata_p0_29__bench,
		n2_odata_p0_30__bench,
		n2_odata_p0_31__bench,
		n2_odata_p0_32__bench,
		n2_odata_p0_33__bench,
		n2_odata_p0_34__bench}),
		.n2_ovalid_p0(n2_ovalid_p0_bench),
		.n3_ordy_p0({n3_ordy_p0_0__bench,
		n3_ordy_p0_1__bench}),
		.n3_odata_p0({n3_odata_p0_0__bench,
		n3_odata_p0_1__bench,
		n3_odata_p0_2__bench,
		n3_odata_p0_3__bench,
		n3_odata_p0_4__bench,
		n3_odata_p0_5__bench,
		n3_odata_p0_6__bench,
		n3_odata_p0_7__bench,
		n3_odata_p0_8__bench,
		n3_odata_p0_9__bench,
		n3_odata_p0_10__bench,
		n3_odata_p0_11__bench,
		n3_odata_p0_12__bench,
		n3_odata_p0_13__bench,
		n3_odata_p0_14__bench,
		n3_odata_p0_15__bench,
		n3_odata_p0_16__bench,
		n3_odata_p0_17__bench,
		n3_odata_p0_18__bench,
		n3_odata_p0_19__bench,
		n3_odata_p0_20__bench,
		n3_odata_p0_21__bench,
		n3_odata_p0_22__bench,
		n3_odata_p0_23__bench,
		n3_odata_p0_24__bench,
		n3_odata_p0_25__bench,
		n3_odata_p0_26__bench,
		n3_odata_p0_27__bench,
		n3_odata_p0_28__bench,
		n3_odata_p0_29__bench,
		n3_odata_p0_30__bench,
		n3_odata_p0_31__bench,
		n3_odata_p0_32__bench,
		n3_odata_p0_33__bench,
		n3_odata_p0_34__bench}),
		.n3_ovalid_p0(n3_ovalid_p0_bench),
		.n4_ordy_p0({n4_ordy_p0_0__bench,
		n4_ordy_p0_1__bench}),
		.n4_odata_p0({n4_odata_p0_0__bench,
		n4_odata_p0_1__bench,
		n4_odata_p0_2__bench,
		n4_odata_p0_3__bench,
		n4_odata_p0_4__bench,
		n4_odata_p0_5__bench,
		n4_odata_p0_6__bench,
		n4_odata_p0_7__bench,
		n4_odata_p0_8__bench,
		n4_odata_p0_9__bench,
		n4_odata_p0_10__bench,
		n4_odata_p0_11__bench,
		n4_odata_p0_12__bench,
		n4_odata_p0_13__bench,
		n4_odata_p0_14__bench,
		n4_odata_p0_15__bench,
		n4_odata_p0_16__bench,
		n4_odata_p0_17__bench,
		n4_odata_p0_18__bench,
		n4_odata_p0_19__bench,
		n4_odata_p0_20__bench,
		n4_odata_p0_21__bench,
		n4_odata_p0_22__bench,
		n4_odata_p0_23__bench,
		n4_odata_p0_24__bench,
		n4_odata_p0_25__bench,
		n4_odata_p0_26__bench,
		n4_odata_p0_27__bench,
		n4_odata_p0_28__bench,
		n4_odata_p0_29__bench,
		n4_odata_p0_30__bench,
		n4_odata_p0_31__bench,
		n4_odata_p0_32__bench,
		n4_odata_p0_33__bench,
		n4_odata_p0_34__bench}),
		.n4_ovalid_p0(n4_ovalid_p0_bench),
		.n5_ordy_p0({n5_ordy_p0_0__bench,
		n5_ordy_p0_1__bench}),
		.n5_odata_p0({n5_odata_p0_0__bench,
		n5_odata_p0_1__bench,
		n5_odata_p0_2__bench,
		n5_odata_p0_3__bench,
		n5_odata_p0_4__bench,
		n5_odata_p0_5__bench,
		n5_odata_p0_6__bench,
		n5_odata_p0_7__bench,
		n5_odata_p0_8__bench,
		n5_odata_p0_9__bench,
		n5_odata_p0_10__bench,
		n5_odata_p0_11__bench,
		n5_odata_p0_12__bench,
		n5_odata_p0_13__bench,
		n5_odata_p0_14__bench,
		n5_odata_p0_15__bench,
		n5_odata_p0_16__bench,
		n5_odata_p0_17__bench,
		n5_odata_p0_18__bench,
		n5_odata_p0_19__bench,
		n5_odata_p0_20__bench,
		n5_odata_p0_21__bench,
		n5_odata_p0_22__bench,
		n5_odata_p0_23__bench,
		n5_odata_p0_24__bench,
		n5_odata_p0_25__bench,
		n5_odata_p0_26__bench,
		n5_odata_p0_27__bench,
		n5_odata_p0_28__bench,
		n5_odata_p0_29__bench,
		n5_odata_p0_30__bench,
		n5_odata_p0_31__bench,
		n5_odata_p0_32__bench,
		n5_odata_p0_33__bench,
		n5_odata_p0_34__bench}),
		.n5_ovalid_p0(n5_ovalid_p0_bench),
		.n6_ordy_p0({n6_ordy_p0_0__bench,
		n6_ordy_p0_1__bench}),
		.n6_odata_p0({n6_odata_p0_0__bench,
		n6_odata_p0_1__bench,
		n6_odata_p0_2__bench,
		n6_odata_p0_3__bench,
		n6_odata_p0_4__bench,
		n6_odata_p0_5__bench,
		n6_odata_p0_6__bench,
		n6_odata_p0_7__bench,
		n6_odata_p0_8__bench,
		n6_odata_p0_9__bench,
		n6_odata_p0_10__bench,
		n6_odata_p0_11__bench,
		n6_odata_p0_12__bench,
		n6_odata_p0_13__bench,
		n6_odata_p0_14__bench,
		n6_odata_p0_15__bench,
		n6_odata_p0_16__bench,
		n6_odata_p0_17__bench,
		n6_odata_p0_18__bench,
		n6_odata_p0_19__bench,
		n6_odata_p0_20__bench,
		n6_odata_p0_21__bench,
		n6_odata_p0_22__bench,
		n6_odata_p0_23__bench,
		n6_odata_p0_24__bench,
		n6_odata_p0_25__bench,
		n6_odata_p0_26__bench,
		n6_odata_p0_27__bench,
		n6_odata_p0_28__bench,
		n6_odata_p0_29__bench,
		n6_odata_p0_30__bench,
		n6_odata_p0_31__bench,
		n6_odata_p0_32__bench,
		n6_odata_p0_33__bench,
		n6_odata_p0_34__bench}),
		.n6_ovalid_p0(n6_ovalid_p0_bench),
		.n7_ordy_p0({n7_ordy_p0_0__bench,
		n7_ordy_p0_1__bench}),
		.n7_odata_p0({n7_odata_p0_0__bench,
		n7_odata_p0_1__bench,
		n7_odata_p0_2__bench,
		n7_odata_p0_3__bench,
		n7_odata_p0_4__bench,
		n7_odata_p0_5__bench,
		n7_odata_p0_6__bench,
		n7_odata_p0_7__bench,
		n7_odata_p0_8__bench,
		n7_odata_p0_9__bench,
		n7_odata_p0_10__bench,
		n7_odata_p0_11__bench,
		n7_odata_p0_12__bench,
		n7_odata_p0_13__bench,
		n7_odata_p0_14__bench,
		n7_odata_p0_15__bench,
		n7_odata_p0_16__bench,
		n7_odata_p0_17__bench,
		n7_odata_p0_18__bench,
		n7_odata_p0_19__bench,
		n7_odata_p0_20__bench,
		n7_odata_p0_21__bench,
		n7_odata_p0_22__bench,
		n7_odata_p0_23__bench,
		n7_odata_p0_24__bench,
		n7_odata_p0_25__bench,
		n7_odata_p0_26__bench,
		n7_odata_p0_27__bench,
		n7_odata_p0_28__bench,
		n7_odata_p0_29__bench,
		n7_odata_p0_30__bench,
		n7_odata_p0_31__bench,
		n7_odata_p0_32__bench,
		n7_odata_p0_33__bench,
		n7_odata_p0_34__bench}),
		.n7_ovalid_p0(n7_ovalid_p0_bench),
		.n8_ordy_p0({n8_ordy_p0_0__bench,
		n8_ordy_p0_1__bench}),
		.n8_odata_p0({n8_odata_p0_0__bench,
		n8_odata_p0_1__bench,
		n8_odata_p0_2__bench,
		n8_odata_p0_3__bench,
		n8_odata_p0_4__bench,
		n8_odata_p0_5__bench,
		n8_odata_p0_6__bench,
		n8_odata_p0_7__bench,
		n8_odata_p0_8__bench,
		n8_odata_p0_9__bench,
		n8_odata_p0_10__bench,
		n8_odata_p0_11__bench,
		n8_odata_p0_12__bench,
		n8_odata_p0_13__bench,
		n8_odata_p0_14__bench,
		n8_odata_p0_15__bench,
		n8_odata_p0_16__bench,
		n8_odata_p0_17__bench,
		n8_odata_p0_18__bench,
		n8_odata_p0_19__bench,
		n8_odata_p0_20__bench,
		n8_odata_p0_21__bench,
		n8_odata_p0_22__bench,
		n8_odata_p0_23__bench,
		n8_odata_p0_24__bench,
		n8_odata_p0_25__bench,
		n8_odata_p0_26__bench,
		n8_odata_p0_27__bench,
		n8_odata_p0_28__bench,
		n8_odata_p0_29__bench,
		n8_odata_p0_30__bench,
		n8_odata_p0_31__bench,
		n8_odata_p0_32__bench,
		n8_odata_p0_33__bench,
		n8_odata_p0_34__bench}),
		.n8_ovalid_p0(n8_ovalid_p0_bench)
	); 
// ----- End reference Benchmark Instanication -------

// ----- Clock 'clk' Initialization -------
	initial begin
		clk[0] <= 1'b0;
		while(1) begin
			#1
			clk[0] <= !clk[0];
		end
	end

// ----- Begin reset signal generation -----
// ----- End reset signal generation -----

// ----- Input Initialization -------
	initial begin
		n0_idata_p0_0_ <= 1'b0;
		n0_idata_p0_1_ <= 1'b0;
		n0_idata_p0_2_ <= 1'b0;
		n0_idata_p0_3_ <= 1'b0;
		n0_idata_p0_4_ <= 1'b0;
		n0_idata_p0_5_ <= 1'b0;
		n0_idata_p0_6_ <= 1'b0;
		n0_idata_p0_7_ <= 1'b0;
		n0_idata_p0_8_ <= 1'b0;
		n0_idata_p0_9_ <= 1'b0;
		n0_idata_p0_10_ <= 1'b0;
		n0_idata_p0_11_ <= 1'b0;
		n0_idata_p0_12_ <= 1'b0;
		n0_idata_p0_13_ <= 1'b0;
		n0_idata_p0_14_ <= 1'b0;
		n0_idata_p0_15_ <= 1'b0;
		n0_idata_p0_16_ <= 1'b0;
		n0_idata_p0_17_ <= 1'b0;
		n0_idata_p0_18_ <= 1'b0;
		n0_idata_p0_19_ <= 1'b0;
		n0_idata_p0_20_ <= 1'b0;
		n0_idata_p0_21_ <= 1'b0;
		n0_idata_p0_22_ <= 1'b0;
		n0_idata_p0_23_ <= 1'b0;
		n0_idata_p0_24_ <= 1'b0;
		n0_idata_p0_25_ <= 1'b0;
		n0_idata_p0_26_ <= 1'b0;
		n0_idata_p0_27_ <= 1'b0;
		n0_idata_p0_28_ <= 1'b0;
		n0_idata_p0_29_ <= 1'b0;
		n0_idata_p0_30_ <= 1'b0;
		n0_idata_p0_31_ <= 1'b0;
		n0_idata_p0_32_ <= 1'b0;
		n0_idata_p0_33_ <= 1'b0;
		n0_idata_p0_34_ <= 1'b0;
		n0_ivalid_p0 <= 1'b0;
		n0_ivch_p0 <= 1'b0;
		n1_idata_p0_0_ <= 1'b0;
		n1_idata_p0_1_ <= 1'b0;
		n1_idata_p0_2_ <= 1'b0;
		n1_idata_p0_3_ <= 1'b0;
		n1_idata_p0_4_ <= 1'b0;
		n1_idata_p0_5_ <= 1'b0;
		n1_idata_p0_6_ <= 1'b0;
		n1_idata_p0_7_ <= 1'b0;
		n1_idata_p0_8_ <= 1'b0;
		n1_idata_p0_9_ <= 1'b0;
		n1_idata_p0_10_ <= 1'b0;
		n1_idata_p0_11_ <= 1'b0;
		n1_idata_p0_12_ <= 1'b0;
		n1_idata_p0_13_ <= 1'b0;
		n1_idata_p0_14_ <= 1'b0;
		n1_idata_p0_15_ <= 1'b0;
		n1_idata_p0_16_ <= 1'b0;
		n1_idata_p0_17_ <= 1'b0;
		n1_idata_p0_18_ <= 1'b0;
		n1_idata_p0_19_ <= 1'b0;
		n1_idata_p0_20_ <= 1'b0;
		n1_idata_p0_21_ <= 1'b0;
		n1_idata_p0_22_ <= 1'b0;
		n1_idata_p0_23_ <= 1'b0;
		n1_idata_p0_24_ <= 1'b0;
		n1_idata_p0_25_ <= 1'b0;
		n1_idata_p0_26_ <= 1'b0;
		n1_idata_p0_27_ <= 1'b0;
		n1_idata_p0_28_ <= 1'b0;
		n1_idata_p0_29_ <= 1'b0;
		n1_idata_p0_30_ <= 1'b0;
		n1_idata_p0_31_ <= 1'b0;
		n1_idata_p0_32_ <= 1'b0;
		n1_idata_p0_33_ <= 1'b0;
		n1_idata_p0_34_ <= 1'b0;
		n1_ivalid_p0 <= 1'b0;
		n1_ivch_p0 <= 1'b0;
		n2_idata_p0_0_ <= 1'b0;
		n2_idata_p0_1_ <= 1'b0;
		n2_idata_p0_2_ <= 1'b0;
		n2_idata_p0_3_ <= 1'b0;
		n2_idata_p0_4_ <= 1'b0;
		n2_idata_p0_5_ <= 1'b0;
		n2_idata_p0_6_ <= 1'b0;
		n2_idata_p0_7_ <= 1'b0;
		n2_idata_p0_8_ <= 1'b0;
		n2_idata_p0_9_ <= 1'b0;
		n2_idata_p0_10_ <= 1'b0;
		n2_idata_p0_11_ <= 1'b0;
		n2_idata_p0_12_ <= 1'b0;
		n2_idata_p0_13_ <= 1'b0;
		n2_idata_p0_14_ <= 1'b0;
		n2_idata_p0_15_ <= 1'b0;
		n2_idata_p0_16_ <= 1'b0;
		n2_idata_p0_17_ <= 1'b0;
		n2_idata_p0_18_ <= 1'b0;
		n2_idata_p0_19_ <= 1'b0;
		n2_idata_p0_20_ <= 1'b0;
		n2_idata_p0_21_ <= 1'b0;
		n2_idata_p0_22_ <= 1'b0;
		n2_idata_p0_23_ <= 1'b0;
		n2_idata_p0_24_ <= 1'b0;
		n2_idata_p0_25_ <= 1'b0;
		n2_idata_p0_26_ <= 1'b0;
		n2_idata_p0_27_ <= 1'b0;
		n2_idata_p0_28_ <= 1'b0;
		n2_idata_p0_29_ <= 1'b0;
		n2_idata_p0_30_ <= 1'b0;
		n2_idata_p0_31_ <= 1'b0;
		n2_idata_p0_32_ <= 1'b0;
		n2_idata_p0_33_ <= 1'b0;
		n2_idata_p0_34_ <= 1'b0;
		n2_ivalid_p0 <= 1'b0;
		n2_ivch_p0 <= 1'b0;
		n3_idata_p0_0_ <= 1'b0;
		n3_idata_p0_1_ <= 1'b0;
		n3_idata_p0_2_ <= 1'b0;
		n3_idata_p0_3_ <= 1'b0;
		n3_idata_p0_4_ <= 1'b0;
		n3_idata_p0_5_ <= 1'b0;
		n3_idata_p0_6_ <= 1'b0;
		n3_idata_p0_7_ <= 1'b0;
		n3_idata_p0_8_ <= 1'b0;
		n3_idata_p0_9_ <= 1'b0;
		n3_idata_p0_10_ <= 1'b0;
		n3_idata_p0_11_ <= 1'b0;
		n3_idata_p0_12_ <= 1'b0;
		n3_idata_p0_13_ <= 1'b0;
		n3_idata_p0_14_ <= 1'b0;
		n3_idata_p0_15_ <= 1'b0;
		n3_idata_p0_16_ <= 1'b0;
		n3_idata_p0_17_ <= 1'b0;
		n3_idata_p0_18_ <= 1'b0;
		n3_idata_p0_19_ <= 1'b0;
		n3_idata_p0_20_ <= 1'b0;
		n3_idata_p0_21_ <= 1'b0;
		n3_idata_p0_22_ <= 1'b0;
		n3_idata_p0_23_ <= 1'b0;
		n3_idata_p0_24_ <= 1'b0;
		n3_idata_p0_25_ <= 1'b0;
		n3_idata_p0_26_ <= 1'b0;
		n3_idata_p0_27_ <= 1'b0;
		n3_idata_p0_28_ <= 1'b0;
		n3_idata_p0_29_ <= 1'b0;
		n3_idata_p0_30_ <= 1'b0;
		n3_idata_p0_31_ <= 1'b0;
		n3_idata_p0_32_ <= 1'b0;
		n3_idata_p0_33_ <= 1'b0;
		n3_idata_p0_34_ <= 1'b0;
		n3_ivalid_p0 <= 1'b0;
		n3_ivch_p0 <= 1'b0;
		n4_idata_p0_0_ <= 1'b0;
		n4_idata_p0_1_ <= 1'b0;
		n4_idata_p0_2_ <= 1'b0;
		n4_idata_p0_3_ <= 1'b0;
		n4_idata_p0_4_ <= 1'b0;
		n4_idata_p0_5_ <= 1'b0;
		n4_idata_p0_6_ <= 1'b0;
		n4_idata_p0_7_ <= 1'b0;
		n4_idata_p0_8_ <= 1'b0;
		n4_idata_p0_9_ <= 1'b0;
		n4_idata_p0_10_ <= 1'b0;
		n4_idata_p0_11_ <= 1'b0;
		n4_idata_p0_12_ <= 1'b0;
		n4_idata_p0_13_ <= 1'b0;
		n4_idata_p0_14_ <= 1'b0;
		n4_idata_p0_15_ <= 1'b0;
		n4_idata_p0_16_ <= 1'b0;
		n4_idata_p0_17_ <= 1'b0;
		n4_idata_p0_18_ <= 1'b0;
		n4_idata_p0_19_ <= 1'b0;
		n4_idata_p0_20_ <= 1'b0;
		n4_idata_p0_21_ <= 1'b0;
		n4_idata_p0_22_ <= 1'b0;
		n4_idata_p0_23_ <= 1'b0;
		n4_idata_p0_24_ <= 1'b0;
		n4_idata_p0_25_ <= 1'b0;
		n4_idata_p0_26_ <= 1'b0;
		n4_idata_p0_27_ <= 1'b0;
		n4_idata_p0_28_ <= 1'b0;
		n4_idata_p0_29_ <= 1'b0;
		n4_idata_p0_30_ <= 1'b0;
		n4_idata_p0_31_ <= 1'b0;
		n4_idata_p0_32_ <= 1'b0;
		n4_idata_p0_33_ <= 1'b0;
		n4_idata_p0_34_ <= 1'b0;
		n4_ivalid_p0 <= 1'b0;
		n4_ivch_p0 <= 1'b0;
		n5_idata_p0_0_ <= 1'b0;
		n5_idata_p0_1_ <= 1'b0;
		n5_idata_p0_2_ <= 1'b0;
		n5_idata_p0_3_ <= 1'b0;
		n5_idata_p0_4_ <= 1'b0;
		n5_idata_p0_5_ <= 1'b0;
		n5_idata_p0_6_ <= 1'b0;
		n5_idata_p0_7_ <= 1'b0;
		n5_idata_p0_8_ <= 1'b0;
		n5_idata_p0_9_ <= 1'b0;
		n5_idata_p0_10_ <= 1'b0;
		n5_idata_p0_11_ <= 1'b0;
		n5_idata_p0_12_ <= 1'b0;
		n5_idata_p0_13_ <= 1'b0;
		n5_idata_p0_14_ <= 1'b0;
		n5_idata_p0_15_ <= 1'b0;
		n5_idata_p0_16_ <= 1'b0;
		n5_idata_p0_17_ <= 1'b0;
		n5_idata_p0_18_ <= 1'b0;
		n5_idata_p0_19_ <= 1'b0;
		n5_idata_p0_20_ <= 1'b0;
		n5_idata_p0_21_ <= 1'b0;
		n5_idata_p0_22_ <= 1'b0;
		n5_idata_p0_23_ <= 1'b0;
		n5_idata_p0_24_ <= 1'b0;
		n5_idata_p0_25_ <= 1'b0;
		n5_idata_p0_26_ <= 1'b0;
		n5_idata_p0_27_ <= 1'b0;
		n5_idata_p0_28_ <= 1'b0;
		n5_idata_p0_29_ <= 1'b0;
		n5_idata_p0_30_ <= 1'b0;
		n5_idata_p0_31_ <= 1'b0;
		n5_idata_p0_32_ <= 1'b0;
		n5_idata_p0_33_ <= 1'b0;
		n5_idata_p0_34_ <= 1'b0;
		n5_ivalid_p0 <= 1'b0;
		n5_ivch_p0 <= 1'b0;
		n6_idata_p0_0_ <= 1'b0;
		n6_idata_p0_1_ <= 1'b0;
		n6_idata_p0_2_ <= 1'b0;
		n6_idata_p0_3_ <= 1'b0;
		n6_idata_p0_4_ <= 1'b0;
		n6_idata_p0_5_ <= 1'b0;
		n6_idata_p0_6_ <= 1'b0;
		n6_idata_p0_7_ <= 1'b0;
		n6_idata_p0_8_ <= 1'b0;
		n6_idata_p0_9_ <= 1'b0;
		n6_idata_p0_10_ <= 1'b0;
		n6_idata_p0_11_ <= 1'b0;
		n6_idata_p0_12_ <= 1'b0;
		n6_idata_p0_13_ <= 1'b0;
		n6_idata_p0_14_ <= 1'b0;
		n6_idata_p0_15_ <= 1'b0;
		n6_idata_p0_16_ <= 1'b0;
		n6_idata_p0_17_ <= 1'b0;
		n6_idata_p0_18_ <= 1'b0;
		n6_idata_p0_19_ <= 1'b0;
		n6_idata_p0_20_ <= 1'b0;
		n6_idata_p0_21_ <= 1'b0;
		n6_idata_p0_22_ <= 1'b0;
		n6_idata_p0_23_ <= 1'b0;
		n6_idata_p0_24_ <= 1'b0;
		n6_idata_p0_25_ <= 1'b0;
		n6_idata_p0_26_ <= 1'b0;
		n6_idata_p0_27_ <= 1'b0;
		n6_idata_p0_28_ <= 1'b0;
		n6_idata_p0_29_ <= 1'b0;
		n6_idata_p0_30_ <= 1'b0;
		n6_idata_p0_31_ <= 1'b0;
		n6_idata_p0_32_ <= 1'b0;
		n6_idata_p0_33_ <= 1'b0;
		n6_idata_p0_34_ <= 1'b0;
		n6_ivalid_p0 <= 1'b0;
		n6_ivch_p0 <= 1'b0;
		n7_idata_p0_0_ <= 1'b0;
		n7_idata_p0_1_ <= 1'b0;
		n7_idata_p0_2_ <= 1'b0;
		n7_idata_p0_3_ <= 1'b0;
		n7_idata_p0_4_ <= 1'b0;
		n7_idata_p0_5_ <= 1'b0;
		n7_idata_p0_6_ <= 1'b0;
		n7_idata_p0_7_ <= 1'b0;
		n7_idata_p0_8_ <= 1'b0;
		n7_idata_p0_9_ <= 1'b0;
		n7_idata_p0_10_ <= 1'b0;
		n7_idata_p0_11_ <= 1'b0;
		n7_idata_p0_12_ <= 1'b0;
		n7_idata_p0_13_ <= 1'b0;
		n7_idata_p0_14_ <= 1'b0;
		n7_idata_p0_15_ <= 1'b0;
		n7_idata_p0_16_ <= 1'b0;
		n7_idata_p0_17_ <= 1'b0;
		n7_idata_p0_18_ <= 1'b0;
		n7_idata_p0_19_ <= 1'b0;
		n7_idata_p0_20_ <= 1'b0;
		n7_idata_p0_21_ <= 1'b0;
		n7_idata_p0_22_ <= 1'b0;
		n7_idata_p0_23_ <= 1'b0;
		n7_idata_p0_24_ <= 1'b0;
		n7_idata_p0_25_ <= 1'b0;
		n7_idata_p0_26_ <= 1'b0;
		n7_idata_p0_27_ <= 1'b0;
		n7_idata_p0_28_ <= 1'b0;
		n7_idata_p0_29_ <= 1'b0;
		n7_idata_p0_30_ <= 1'b0;
		n7_idata_p0_31_ <= 1'b0;
		n7_idata_p0_32_ <= 1'b0;
		n7_idata_p0_33_ <= 1'b0;
		n7_idata_p0_34_ <= 1'b0;
		n7_ivalid_p0 <= 1'b0;
		n7_ivch_p0 <= 1'b0;
		n8_idata_p0_0_ <= 1'b0;
		n8_idata_p0_1_ <= 1'b0;
		n8_idata_p0_2_ <= 1'b0;
		n8_idata_p0_3_ <= 1'b0;
		n8_idata_p0_4_ <= 1'b0;
		n8_idata_p0_5_ <= 1'b0;
		n8_idata_p0_6_ <= 1'b0;
		n8_idata_p0_7_ <= 1'b0;
		n8_idata_p0_8_ <= 1'b0;
		n8_idata_p0_9_ <= 1'b0;
		n8_idata_p0_10_ <= 1'b0;
		n8_idata_p0_11_ <= 1'b0;
		n8_idata_p0_12_ <= 1'b0;
		n8_idata_p0_13_ <= 1'b0;
		n8_idata_p0_14_ <= 1'b0;
		n8_idata_p0_15_ <= 1'b0;
		n8_idata_p0_16_ <= 1'b0;
		n8_idata_p0_17_ <= 1'b0;
		n8_idata_p0_18_ <= 1'b0;
		n8_idata_p0_19_ <= 1'b0;
		n8_idata_p0_20_ <= 1'b0;
		n8_idata_p0_21_ <= 1'b0;
		n8_idata_p0_22_ <= 1'b0;
		n8_idata_p0_23_ <= 1'b0;
		n8_idata_p0_24_ <= 1'b0;
		n8_idata_p0_25_ <= 1'b0;
		n8_idata_p0_26_ <= 1'b0;
		n8_idata_p0_27_ <= 1'b0;
		n8_idata_p0_28_ <= 1'b0;
		n8_idata_p0_29_ <= 1'b0;
		n8_idata_p0_30_ <= 1'b0;
		n8_idata_p0_31_ <= 1'b0;
		n8_idata_p0_32_ <= 1'b0;
		n8_idata_p0_33_ <= 1'b0;
		n8_idata_p0_34_ <= 1'b0;
		n8_ivalid_p0 <= 1'b0;
		n8_ivch_p0 <= 1'b0;
		rst_ <= 1'b0;

		n0_ordy_p0_0__flag[0] <= 1'b0;
		n0_ordy_p0_1__flag[0] <= 1'b0;
		n0_odata_p0_0__flag[0] <= 1'b0;
		n0_odata_p0_1__flag[0] <= 1'b0;
		n0_odata_p0_2__flag[0] <= 1'b0;
		n0_odata_p0_3__flag[0] <= 1'b0;
		n0_odata_p0_4__flag[0] <= 1'b0;
		n0_odata_p0_5__flag[0] <= 1'b0;
		n0_odata_p0_6__flag[0] <= 1'b0;
		n0_odata_p0_7__flag[0] <= 1'b0;
		n0_odata_p0_8__flag[0] <= 1'b0;
		n0_odata_p0_9__flag[0] <= 1'b0;
		n0_odata_p0_10__flag[0] <= 1'b0;
		n0_odata_p0_11__flag[0] <= 1'b0;
		n0_odata_p0_12__flag[0] <= 1'b0;
		n0_odata_p0_13__flag[0] <= 1'b0;
		n0_odata_p0_14__flag[0] <= 1'b0;
		n0_odata_p0_15__flag[0] <= 1'b0;
		n0_odata_p0_16__flag[0] <= 1'b0;
		n0_odata_p0_17__flag[0] <= 1'b0;
		n0_odata_p0_18__flag[0] <= 1'b0;
		n0_odata_p0_19__flag[0] <= 1'b0;
		n0_odata_p0_20__flag[0] <= 1'b0;
		n0_odata_p0_21__flag[0] <= 1'b0;
		n0_odata_p0_22__flag[0] <= 1'b0;
		n0_odata_p0_23__flag[0] <= 1'b0;
		n0_odata_p0_24__flag[0] <= 1'b0;
		n0_odata_p0_25__flag[0] <= 1'b0;
		n0_odata_p0_26__flag[0] <= 1'b0;
		n0_odata_p0_27__flag[0] <= 1'b0;
		n0_odata_p0_28__flag[0] <= 1'b0;
		n0_odata_p0_29__flag[0] <= 1'b0;
		n0_odata_p0_30__flag[0] <= 1'b0;
		n0_odata_p0_31__flag[0] <= 1'b0;
		n0_odata_p0_32__flag[0] <= 1'b0;
		n0_odata_p0_33__flag[0] <= 1'b0;
		n0_odata_p0_34__flag[0] <= 1'b0;
		n0_ovalid_p0_flag[0] <= 1'b0;
		n1_ordy_p0_0__flag[0] <= 1'b0;
		n1_ordy_p0_1__flag[0] <= 1'b0;
		n1_odata_p0_0__flag[0] <= 1'b0;
		n1_odata_p0_1__flag[0] <= 1'b0;
		n1_odata_p0_2__flag[0] <= 1'b0;
		n1_odata_p0_3__flag[0] <= 1'b0;
		n1_odata_p0_4__flag[0] <= 1'b0;
		n1_odata_p0_5__flag[0] <= 1'b0;
		n1_odata_p0_6__flag[0] <= 1'b0;
		n1_odata_p0_7__flag[0] <= 1'b0;
		n1_odata_p0_8__flag[0] <= 1'b0;
		n1_odata_p0_9__flag[0] <= 1'b0;
		n1_odata_p0_10__flag[0] <= 1'b0;
		n1_odata_p0_11__flag[0] <= 1'b0;
		n1_odata_p0_12__flag[0] <= 1'b0;
		n1_odata_p0_13__flag[0] <= 1'b0;
		n1_odata_p0_14__flag[0] <= 1'b0;
		n1_odata_p0_15__flag[0] <= 1'b0;
		n1_odata_p0_16__flag[0] <= 1'b0;
		n1_odata_p0_17__flag[0] <= 1'b0;
		n1_odata_p0_18__flag[0] <= 1'b0;
		n1_odata_p0_19__flag[0] <= 1'b0;
		n1_odata_p0_20__flag[0] <= 1'b0;
		n1_odata_p0_21__flag[0] <= 1'b0;
		n1_odata_p0_22__flag[0] <= 1'b0;
		n1_odata_p0_23__flag[0] <= 1'b0;
		n1_odata_p0_24__flag[0] <= 1'b0;
		n1_odata_p0_25__flag[0] <= 1'b0;
		n1_odata_p0_26__flag[0] <= 1'b0;
		n1_odata_p0_27__flag[0] <= 1'b0;
		n1_odata_p0_28__flag[0] <= 1'b0;
		n1_odata_p0_29__flag[0] <= 1'b0;
		n1_odata_p0_30__flag[0] <= 1'b0;
		n1_odata_p0_31__flag[0] <= 1'b0;
		n1_odata_p0_32__flag[0] <= 1'b0;
		n1_odata_p0_33__flag[0] <= 1'b0;
		n1_odata_p0_34__flag[0] <= 1'b0;
		n1_ovalid_p0_flag[0] <= 1'b0;
		n2_ordy_p0_0__flag[0] <= 1'b0;
		n2_ordy_p0_1__flag[0] <= 1'b0;
		n2_odata_p0_0__flag[0] <= 1'b0;
		n2_odata_p0_1__flag[0] <= 1'b0;
		n2_odata_p0_2__flag[0] <= 1'b0;
		n2_odata_p0_3__flag[0] <= 1'b0;
		n2_odata_p0_4__flag[0] <= 1'b0;
		n2_odata_p0_5__flag[0] <= 1'b0;
		n2_odata_p0_6__flag[0] <= 1'b0;
		n2_odata_p0_7__flag[0] <= 1'b0;
		n2_odata_p0_8__flag[0] <= 1'b0;
		n2_odata_p0_9__flag[0] <= 1'b0;
		n2_odata_p0_10__flag[0] <= 1'b0;
		n2_odata_p0_11__flag[0] <= 1'b0;
		n2_odata_p0_12__flag[0] <= 1'b0;
		n2_odata_p0_13__flag[0] <= 1'b0;
		n2_odata_p0_14__flag[0] <= 1'b0;
		n2_odata_p0_15__flag[0] <= 1'b0;
		n2_odata_p0_16__flag[0] <= 1'b0;
		n2_odata_p0_17__flag[0] <= 1'b0;
		n2_odata_p0_18__flag[0] <= 1'b0;
		n2_odata_p0_19__flag[0] <= 1'b0;
		n2_odata_p0_20__flag[0] <= 1'b0;
		n2_odata_p0_21__flag[0] <= 1'b0;
		n2_odata_p0_22__flag[0] <= 1'b0;
		n2_odata_p0_23__flag[0] <= 1'b0;
		n2_odata_p0_24__flag[0] <= 1'b0;
		n2_odata_p0_25__flag[0] <= 1'b0;
		n2_odata_p0_26__flag[0] <= 1'b0;
		n2_odata_p0_27__flag[0] <= 1'b0;
		n2_odata_p0_28__flag[0] <= 1'b0;
		n2_odata_p0_29__flag[0] <= 1'b0;
		n2_odata_p0_30__flag[0] <= 1'b0;
		n2_odata_p0_31__flag[0] <= 1'b0;
		n2_odata_p0_32__flag[0] <= 1'b0;
		n2_odata_p0_33__flag[0] <= 1'b0;
		n2_odata_p0_34__flag[0] <= 1'b0;
		n2_ovalid_p0_flag[0] <= 1'b0;
		n3_ordy_p0_0__flag[0] <= 1'b0;
		n3_ordy_p0_1__flag[0] <= 1'b0;
		n3_odata_p0_0__flag[0] <= 1'b0;
		n3_odata_p0_1__flag[0] <= 1'b0;
		n3_odata_p0_2__flag[0] <= 1'b0;
		n3_odata_p0_3__flag[0] <= 1'b0;
		n3_odata_p0_4__flag[0] <= 1'b0;
		n3_odata_p0_5__flag[0] <= 1'b0;
		n3_odata_p0_6__flag[0] <= 1'b0;
		n3_odata_p0_7__flag[0] <= 1'b0;
		n3_odata_p0_8__flag[0] <= 1'b0;
		n3_odata_p0_9__flag[0] <= 1'b0;
		n3_odata_p0_10__flag[0] <= 1'b0;
		n3_odata_p0_11__flag[0] <= 1'b0;
		n3_odata_p0_12__flag[0] <= 1'b0;
		n3_odata_p0_13__flag[0] <= 1'b0;
		n3_odata_p0_14__flag[0] <= 1'b0;
		n3_odata_p0_15__flag[0] <= 1'b0;
		n3_odata_p0_16__flag[0] <= 1'b0;
		n3_odata_p0_17__flag[0] <= 1'b0;
		n3_odata_p0_18__flag[0] <= 1'b0;
		n3_odata_p0_19__flag[0] <= 1'b0;
		n3_odata_p0_20__flag[0] <= 1'b0;
		n3_odata_p0_21__flag[0] <= 1'b0;
		n3_odata_p0_22__flag[0] <= 1'b0;
		n3_odata_p0_23__flag[0] <= 1'b0;
		n3_odata_p0_24__flag[0] <= 1'b0;
		n3_odata_p0_25__flag[0] <= 1'b0;
		n3_odata_p0_26__flag[0] <= 1'b0;
		n3_odata_p0_27__flag[0] <= 1'b0;
		n3_odata_p0_28__flag[0] <= 1'b0;
		n3_odata_p0_29__flag[0] <= 1'b0;
		n3_odata_p0_30__flag[0] <= 1'b0;
		n3_odata_p0_31__flag[0] <= 1'b0;
		n3_odata_p0_32__flag[0] <= 1'b0;
		n3_odata_p0_33__flag[0] <= 1'b0;
		n3_odata_p0_34__flag[0] <= 1'b0;
		n3_ovalid_p0_flag[0] <= 1'b0;
		n4_ordy_p0_0__flag[0] <= 1'b0;
		n4_ordy_p0_1__flag[0] <= 1'b0;
		n4_odata_p0_0__flag[0] <= 1'b0;
		n4_odata_p0_1__flag[0] <= 1'b0;
		n4_odata_p0_2__flag[0] <= 1'b0;
		n4_odata_p0_3__flag[0] <= 1'b0;
		n4_odata_p0_4__flag[0] <= 1'b0;
		n4_odata_p0_5__flag[0] <= 1'b0;
		n4_odata_p0_6__flag[0] <= 1'b0;
		n4_odata_p0_7__flag[0] <= 1'b0;
		n4_odata_p0_8__flag[0] <= 1'b0;
		n4_odata_p0_9__flag[0] <= 1'b0;
		n4_odata_p0_10__flag[0] <= 1'b0;
		n4_odata_p0_11__flag[0] <= 1'b0;
		n4_odata_p0_12__flag[0] <= 1'b0;
		n4_odata_p0_13__flag[0] <= 1'b0;
		n4_odata_p0_14__flag[0] <= 1'b0;
		n4_odata_p0_15__flag[0] <= 1'b0;
		n4_odata_p0_16__flag[0] <= 1'b0;
		n4_odata_p0_17__flag[0] <= 1'b0;
		n4_odata_p0_18__flag[0] <= 1'b0;
		n4_odata_p0_19__flag[0] <= 1'b0;
		n4_odata_p0_20__flag[0] <= 1'b0;
		n4_odata_p0_21__flag[0] <= 1'b0;
		n4_odata_p0_22__flag[0] <= 1'b0;
		n4_odata_p0_23__flag[0] <= 1'b0;
		n4_odata_p0_24__flag[0] <= 1'b0;
		n4_odata_p0_25__flag[0] <= 1'b0;
		n4_odata_p0_26__flag[0] <= 1'b0;
		n4_odata_p0_27__flag[0] <= 1'b0;
		n4_odata_p0_28__flag[0] <= 1'b0;
		n4_odata_p0_29__flag[0] <= 1'b0;
		n4_odata_p0_30__flag[0] <= 1'b0;
		n4_odata_p0_31__flag[0] <= 1'b0;
		n4_odata_p0_32__flag[0] <= 1'b0;
		n4_odata_p0_33__flag[0] <= 1'b0;
		n4_odata_p0_34__flag[0] <= 1'b0;
		n4_ovalid_p0_flag[0] <= 1'b0;
		n5_ordy_p0_0__flag[0] <= 1'b0;
		n5_ordy_p0_1__flag[0] <= 1'b0;
		n5_odata_p0_0__flag[0] <= 1'b0;
		n5_odata_p0_1__flag[0] <= 1'b0;
		n5_odata_p0_2__flag[0] <= 1'b0;
		n5_odata_p0_3__flag[0] <= 1'b0;
		n5_odata_p0_4__flag[0] <= 1'b0;
		n5_odata_p0_5__flag[0] <= 1'b0;
		n5_odata_p0_6__flag[0] <= 1'b0;
		n5_odata_p0_7__flag[0] <= 1'b0;
		n5_odata_p0_8__flag[0] <= 1'b0;
		n5_odata_p0_9__flag[0] <= 1'b0;
		n5_odata_p0_10__flag[0] <= 1'b0;
		n5_odata_p0_11__flag[0] <= 1'b0;
		n5_odata_p0_12__flag[0] <= 1'b0;
		n5_odata_p0_13__flag[0] <= 1'b0;
		n5_odata_p0_14__flag[0] <= 1'b0;
		n5_odata_p0_15__flag[0] <= 1'b0;
		n5_odata_p0_16__flag[0] <= 1'b0;
		n5_odata_p0_17__flag[0] <= 1'b0;
		n5_odata_p0_18__flag[0] <= 1'b0;
		n5_odata_p0_19__flag[0] <= 1'b0;
		n5_odata_p0_20__flag[0] <= 1'b0;
		n5_odata_p0_21__flag[0] <= 1'b0;
		n5_odata_p0_22__flag[0] <= 1'b0;
		n5_odata_p0_23__flag[0] <= 1'b0;
		n5_odata_p0_24__flag[0] <= 1'b0;
		n5_odata_p0_25__flag[0] <= 1'b0;
		n5_odata_p0_26__flag[0] <= 1'b0;
		n5_odata_p0_27__flag[0] <= 1'b0;
		n5_odata_p0_28__flag[0] <= 1'b0;
		n5_odata_p0_29__flag[0] <= 1'b0;
		n5_odata_p0_30__flag[0] <= 1'b0;
		n5_odata_p0_31__flag[0] <= 1'b0;
		n5_odata_p0_32__flag[0] <= 1'b0;
		n5_odata_p0_33__flag[0] <= 1'b0;
		n5_odata_p0_34__flag[0] <= 1'b0;
		n5_ovalid_p0_flag[0] <= 1'b0;
		n6_ordy_p0_0__flag[0] <= 1'b0;
		n6_ordy_p0_1__flag[0] <= 1'b0;
		n6_odata_p0_0__flag[0] <= 1'b0;
		n6_odata_p0_1__flag[0] <= 1'b0;
		n6_odata_p0_2__flag[0] <= 1'b0;
		n6_odata_p0_3__flag[0] <= 1'b0;
		n6_odata_p0_4__flag[0] <= 1'b0;
		n6_odata_p0_5__flag[0] <= 1'b0;
		n6_odata_p0_6__flag[0] <= 1'b0;
		n6_odata_p0_7__flag[0] <= 1'b0;
		n6_odata_p0_8__flag[0] <= 1'b0;
		n6_odata_p0_9__flag[0] <= 1'b0;
		n6_odata_p0_10__flag[0] <= 1'b0;
		n6_odata_p0_11__flag[0] <= 1'b0;
		n6_odata_p0_12__flag[0] <= 1'b0;
		n6_odata_p0_13__flag[0] <= 1'b0;
		n6_odata_p0_14__flag[0] <= 1'b0;
		n6_odata_p0_15__flag[0] <= 1'b0;
		n6_odata_p0_16__flag[0] <= 1'b0;
		n6_odata_p0_17__flag[0] <= 1'b0;
		n6_odata_p0_18__flag[0] <= 1'b0;
		n6_odata_p0_19__flag[0] <= 1'b0;
		n6_odata_p0_20__flag[0] <= 1'b0;
		n6_odata_p0_21__flag[0] <= 1'b0;
		n6_odata_p0_22__flag[0] <= 1'b0;
		n6_odata_p0_23__flag[0] <= 1'b0;
		n6_odata_p0_24__flag[0] <= 1'b0;
		n6_odata_p0_25__flag[0] <= 1'b0;
		n6_odata_p0_26__flag[0] <= 1'b0;
		n6_odata_p0_27__flag[0] <= 1'b0;
		n6_odata_p0_28__flag[0] <= 1'b0;
		n6_odata_p0_29__flag[0] <= 1'b0;
		n6_odata_p0_30__flag[0] <= 1'b0;
		n6_odata_p0_31__flag[0] <= 1'b0;
		n6_odata_p0_32__flag[0] <= 1'b0;
		n6_odata_p0_33__flag[0] <= 1'b0;
		n6_odata_p0_34__flag[0] <= 1'b0;
		n6_ovalid_p0_flag[0] <= 1'b0;
		n7_ordy_p0_0__flag[0] <= 1'b0;
		n7_ordy_p0_1__flag[0] <= 1'b0;
		n7_odata_p0_0__flag[0] <= 1'b0;
		n7_odata_p0_1__flag[0] <= 1'b0;
		n7_odata_p0_2__flag[0] <= 1'b0;
		n7_odata_p0_3__flag[0] <= 1'b0;
		n7_odata_p0_4__flag[0] <= 1'b0;
		n7_odata_p0_5__flag[0] <= 1'b0;
		n7_odata_p0_6__flag[0] <= 1'b0;
		n7_odata_p0_7__flag[0] <= 1'b0;
		n7_odata_p0_8__flag[0] <= 1'b0;
		n7_odata_p0_9__flag[0] <= 1'b0;
		n7_odata_p0_10__flag[0] <= 1'b0;
		n7_odata_p0_11__flag[0] <= 1'b0;
		n7_odata_p0_12__flag[0] <= 1'b0;
		n7_odata_p0_13__flag[0] <= 1'b0;
		n7_odata_p0_14__flag[0] <= 1'b0;
		n7_odata_p0_15__flag[0] <= 1'b0;
		n7_odata_p0_16__flag[0] <= 1'b0;
		n7_odata_p0_17__flag[0] <= 1'b0;
		n7_odata_p0_18__flag[0] <= 1'b0;
		n7_odata_p0_19__flag[0] <= 1'b0;
		n7_odata_p0_20__flag[0] <= 1'b0;
		n7_odata_p0_21__flag[0] <= 1'b0;
		n7_odata_p0_22__flag[0] <= 1'b0;
		n7_odata_p0_23__flag[0] <= 1'b0;
		n7_odata_p0_24__flag[0] <= 1'b0;
		n7_odata_p0_25__flag[0] <= 1'b0;
		n7_odata_p0_26__flag[0] <= 1'b0;
		n7_odata_p0_27__flag[0] <= 1'b0;
		n7_odata_p0_28__flag[0] <= 1'b0;
		n7_odata_p0_29__flag[0] <= 1'b0;
		n7_odata_p0_30__flag[0] <= 1'b0;
		n7_odata_p0_31__flag[0] <= 1'b0;
		n7_odata_p0_32__flag[0] <= 1'b0;
		n7_odata_p0_33__flag[0] <= 1'b0;
		n7_odata_p0_34__flag[0] <= 1'b0;
		n7_ovalid_p0_flag[0] <= 1'b0;
		n8_ordy_p0_0__flag[0] <= 1'b0;
		n8_ordy_p0_1__flag[0] <= 1'b0;
		n8_odata_p0_0__flag[0] <= 1'b0;
		n8_odata_p0_1__flag[0] <= 1'b0;
		n8_odata_p0_2__flag[0] <= 1'b0;
		n8_odata_p0_3__flag[0] <= 1'b0;
		n8_odata_p0_4__flag[0] <= 1'b0;
		n8_odata_p0_5__flag[0] <= 1'b0;
		n8_odata_p0_6__flag[0] <= 1'b0;
		n8_odata_p0_7__flag[0] <= 1'b0;
		n8_odata_p0_8__flag[0] <= 1'b0;
		n8_odata_p0_9__flag[0] <= 1'b0;
		n8_odata_p0_10__flag[0] <= 1'b0;
		n8_odata_p0_11__flag[0] <= 1'b0;
		n8_odata_p0_12__flag[0] <= 1'b0;
		n8_odata_p0_13__flag[0] <= 1'b0;
		n8_odata_p0_14__flag[0] <= 1'b0;
		n8_odata_p0_15__flag[0] <= 1'b0;
		n8_odata_p0_16__flag[0] <= 1'b0;
		n8_odata_p0_17__flag[0] <= 1'b0;
		n8_odata_p0_18__flag[0] <= 1'b0;
		n8_odata_p0_19__flag[0] <= 1'b0;
		n8_odata_p0_20__flag[0] <= 1'b0;
		n8_odata_p0_21__flag[0] <= 1'b0;
		n8_odata_p0_22__flag[0] <= 1'b0;
		n8_odata_p0_23__flag[0] <= 1'b0;
		n8_odata_p0_24__flag[0] <= 1'b0;
		n8_odata_p0_25__flag[0] <= 1'b0;
		n8_odata_p0_26__flag[0] <= 1'b0;
		n8_odata_p0_27__flag[0] <= 1'b0;
		n8_odata_p0_28__flag[0] <= 1'b0;
		n8_odata_p0_29__flag[0] <= 1'b0;
		n8_odata_p0_30__flag[0] <= 1'b0;
		n8_odata_p0_31__flag[0] <= 1'b0;
		n8_odata_p0_32__flag[0] <= 1'b0;
		n8_odata_p0_33__flag[0] <= 1'b0;
		n8_odata_p0_34__flag[0] <= 1'b0;
		n8_ovalid_p0_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge clk[0]) begin
		n0_idata_p0_0_ <= $random;
		n0_idata_p0_1_ <= $random;
		n0_idata_p0_2_ <= $random;
		n0_idata_p0_3_ <= $random;
		n0_idata_p0_4_ <= $random;
		n0_idata_p0_5_ <= $random;
		n0_idata_p0_6_ <= $random;
		n0_idata_p0_7_ <= $random;
		n0_idata_p0_8_ <= $random;
		n0_idata_p0_9_ <= $random;
		n0_idata_p0_10_ <= $random;
		n0_idata_p0_11_ <= $random;
		n0_idata_p0_12_ <= $random;
		n0_idata_p0_13_ <= $random;
		n0_idata_p0_14_ <= $random;
		n0_idata_p0_15_ <= $random;
		n0_idata_p0_16_ <= $random;
		n0_idata_p0_17_ <= $random;
		n0_idata_p0_18_ <= $random;
		n0_idata_p0_19_ <= $random;
		n0_idata_p0_20_ <= $random;
		n0_idata_p0_21_ <= $random;
		n0_idata_p0_22_ <= $random;
		n0_idata_p0_23_ <= $random;
		n0_idata_p0_24_ <= $random;
		n0_idata_p0_25_ <= $random;
		n0_idata_p0_26_ <= $random;
		n0_idata_p0_27_ <= $random;
		n0_idata_p0_28_ <= $random;
		n0_idata_p0_29_ <= $random;
		n0_idata_p0_30_ <= $random;
		n0_idata_p0_31_ <= $random;
		n0_idata_p0_32_ <= $random;
		n0_idata_p0_33_ <= $random;
		n0_idata_p0_34_ <= $random;
		n0_ivalid_p0 <= $random;
		n0_ivch_p0 <= $random;
		n1_idata_p0_0_ <= $random;
		n1_idata_p0_1_ <= $random;
		n1_idata_p0_2_ <= $random;
		n1_idata_p0_3_ <= $random;
		n1_idata_p0_4_ <= $random;
		n1_idata_p0_5_ <= $random;
		n1_idata_p0_6_ <= $random;
		n1_idata_p0_7_ <= $random;
		n1_idata_p0_8_ <= $random;
		n1_idata_p0_9_ <= $random;
		n1_idata_p0_10_ <= $random;
		n1_idata_p0_11_ <= $random;
		n1_idata_p0_12_ <= $random;
		n1_idata_p0_13_ <= $random;
		n1_idata_p0_14_ <= $random;
		n1_idata_p0_15_ <= $random;
		n1_idata_p0_16_ <= $random;
		n1_idata_p0_17_ <= $random;
		n1_idata_p0_18_ <= $random;
		n1_idata_p0_19_ <= $random;
		n1_idata_p0_20_ <= $random;
		n1_idata_p0_21_ <= $random;
		n1_idata_p0_22_ <= $random;
		n1_idata_p0_23_ <= $random;
		n1_idata_p0_24_ <= $random;
		n1_idata_p0_25_ <= $random;
		n1_idata_p0_26_ <= $random;
		n1_idata_p0_27_ <= $random;
		n1_idata_p0_28_ <= $random;
		n1_idata_p0_29_ <= $random;
		n1_idata_p0_30_ <= $random;
		n1_idata_p0_31_ <= $random;
		n1_idata_p0_32_ <= $random;
		n1_idata_p0_33_ <= $random;
		n1_idata_p0_34_ <= $random;
		n1_ivalid_p0 <= $random;
		n1_ivch_p0 <= $random;
		n2_idata_p0_0_ <= $random;
		n2_idata_p0_1_ <= $random;
		n2_idata_p0_2_ <= $random;
		n2_idata_p0_3_ <= $random;
		n2_idata_p0_4_ <= $random;
		n2_idata_p0_5_ <= $random;
		n2_idata_p0_6_ <= $random;
		n2_idata_p0_7_ <= $random;
		n2_idata_p0_8_ <= $random;
		n2_idata_p0_9_ <= $random;
		n2_idata_p0_10_ <= $random;
		n2_idata_p0_11_ <= $random;
		n2_idata_p0_12_ <= $random;
		n2_idata_p0_13_ <= $random;
		n2_idata_p0_14_ <= $random;
		n2_idata_p0_15_ <= $random;
		n2_idata_p0_16_ <= $random;
		n2_idata_p0_17_ <= $random;
		n2_idata_p0_18_ <= $random;
		n2_idata_p0_19_ <= $random;
		n2_idata_p0_20_ <= $random;
		n2_idata_p0_21_ <= $random;
		n2_idata_p0_22_ <= $random;
		n2_idata_p0_23_ <= $random;
		n2_idata_p0_24_ <= $random;
		n2_idata_p0_25_ <= $random;
		n2_idata_p0_26_ <= $random;
		n2_idata_p0_27_ <= $random;
		n2_idata_p0_28_ <= $random;
		n2_idata_p0_29_ <= $random;
		n2_idata_p0_30_ <= $random;
		n2_idata_p0_31_ <= $random;
		n2_idata_p0_32_ <= $random;
		n2_idata_p0_33_ <= $random;
		n2_idata_p0_34_ <= $random;
		n2_ivalid_p0 <= $random;
		n2_ivch_p0 <= $random;
		n3_idata_p0_0_ <= $random;
		n3_idata_p0_1_ <= $random;
		n3_idata_p0_2_ <= $random;
		n3_idata_p0_3_ <= $random;
		n3_idata_p0_4_ <= $random;
		n3_idata_p0_5_ <= $random;
		n3_idata_p0_6_ <= $random;
		n3_idata_p0_7_ <= $random;
		n3_idata_p0_8_ <= $random;
		n3_idata_p0_9_ <= $random;
		n3_idata_p0_10_ <= $random;
		n3_idata_p0_11_ <= $random;
		n3_idata_p0_12_ <= $random;
		n3_idata_p0_13_ <= $random;
		n3_idata_p0_14_ <= $random;
		n3_idata_p0_15_ <= $random;
		n3_idata_p0_16_ <= $random;
		n3_idata_p0_17_ <= $random;
		n3_idata_p0_18_ <= $random;
		n3_idata_p0_19_ <= $random;
		n3_idata_p0_20_ <= $random;
		n3_idata_p0_21_ <= $random;
		n3_idata_p0_22_ <= $random;
		n3_idata_p0_23_ <= $random;
		n3_idata_p0_24_ <= $random;
		n3_idata_p0_25_ <= $random;
		n3_idata_p0_26_ <= $random;
		n3_idata_p0_27_ <= $random;
		n3_idata_p0_28_ <= $random;
		n3_idata_p0_29_ <= $random;
		n3_idata_p0_30_ <= $random;
		n3_idata_p0_31_ <= $random;
		n3_idata_p0_32_ <= $random;
		n3_idata_p0_33_ <= $random;
		n3_idata_p0_34_ <= $random;
		n3_ivalid_p0 <= $random;
		n3_ivch_p0 <= $random;
		n4_idata_p0_0_ <= $random;
		n4_idata_p0_1_ <= $random;
		n4_idata_p0_2_ <= $random;
		n4_idata_p0_3_ <= $random;
		n4_idata_p0_4_ <= $random;
		n4_idata_p0_5_ <= $random;
		n4_idata_p0_6_ <= $random;
		n4_idata_p0_7_ <= $random;
		n4_idata_p0_8_ <= $random;
		n4_idata_p0_9_ <= $random;
		n4_idata_p0_10_ <= $random;
		n4_idata_p0_11_ <= $random;
		n4_idata_p0_12_ <= $random;
		n4_idata_p0_13_ <= $random;
		n4_idata_p0_14_ <= $random;
		n4_idata_p0_15_ <= $random;
		n4_idata_p0_16_ <= $random;
		n4_idata_p0_17_ <= $random;
		n4_idata_p0_18_ <= $random;
		n4_idata_p0_19_ <= $random;
		n4_idata_p0_20_ <= $random;
		n4_idata_p0_21_ <= $random;
		n4_idata_p0_22_ <= $random;
		n4_idata_p0_23_ <= $random;
		n4_idata_p0_24_ <= $random;
		n4_idata_p0_25_ <= $random;
		n4_idata_p0_26_ <= $random;
		n4_idata_p0_27_ <= $random;
		n4_idata_p0_28_ <= $random;
		n4_idata_p0_29_ <= $random;
		n4_idata_p0_30_ <= $random;
		n4_idata_p0_31_ <= $random;
		n4_idata_p0_32_ <= $random;
		n4_idata_p0_33_ <= $random;
		n4_idata_p0_34_ <= $random;
		n4_ivalid_p0 <= $random;
		n4_ivch_p0 <= $random;
		n5_idata_p0_0_ <= $random;
		n5_idata_p0_1_ <= $random;
		n5_idata_p0_2_ <= $random;
		n5_idata_p0_3_ <= $random;
		n5_idata_p0_4_ <= $random;
		n5_idata_p0_5_ <= $random;
		n5_idata_p0_6_ <= $random;
		n5_idata_p0_7_ <= $random;
		n5_idata_p0_8_ <= $random;
		n5_idata_p0_9_ <= $random;
		n5_idata_p0_10_ <= $random;
		n5_idata_p0_11_ <= $random;
		n5_idata_p0_12_ <= $random;
		n5_idata_p0_13_ <= $random;
		n5_idata_p0_14_ <= $random;
		n5_idata_p0_15_ <= $random;
		n5_idata_p0_16_ <= $random;
		n5_idata_p0_17_ <= $random;
		n5_idata_p0_18_ <= $random;
		n5_idata_p0_19_ <= $random;
		n5_idata_p0_20_ <= $random;
		n5_idata_p0_21_ <= $random;
		n5_idata_p0_22_ <= $random;
		n5_idata_p0_23_ <= $random;
		n5_idata_p0_24_ <= $random;
		n5_idata_p0_25_ <= $random;
		n5_idata_p0_26_ <= $random;
		n5_idata_p0_27_ <= $random;
		n5_idata_p0_28_ <= $random;
		n5_idata_p0_29_ <= $random;
		n5_idata_p0_30_ <= $random;
		n5_idata_p0_31_ <= $random;
		n5_idata_p0_32_ <= $random;
		n5_idata_p0_33_ <= $random;
		n5_idata_p0_34_ <= $random;
		n5_ivalid_p0 <= $random;
		n5_ivch_p0 <= $random;
		n6_idata_p0_0_ <= $random;
		n6_idata_p0_1_ <= $random;
		n6_idata_p0_2_ <= $random;
		n6_idata_p0_3_ <= $random;
		n6_idata_p0_4_ <= $random;
		n6_idata_p0_5_ <= $random;
		n6_idata_p0_6_ <= $random;
		n6_idata_p0_7_ <= $random;
		n6_idata_p0_8_ <= $random;
		n6_idata_p0_9_ <= $random;
		n6_idata_p0_10_ <= $random;
		n6_idata_p0_11_ <= $random;
		n6_idata_p0_12_ <= $random;
		n6_idata_p0_13_ <= $random;
		n6_idata_p0_14_ <= $random;
		n6_idata_p0_15_ <= $random;
		n6_idata_p0_16_ <= $random;
		n6_idata_p0_17_ <= $random;
		n6_idata_p0_18_ <= $random;
		n6_idata_p0_19_ <= $random;
		n6_idata_p0_20_ <= $random;
		n6_idata_p0_21_ <= $random;
		n6_idata_p0_22_ <= $random;
		n6_idata_p0_23_ <= $random;
		n6_idata_p0_24_ <= $random;
		n6_idata_p0_25_ <= $random;
		n6_idata_p0_26_ <= $random;
		n6_idata_p0_27_ <= $random;
		n6_idata_p0_28_ <= $random;
		n6_idata_p0_29_ <= $random;
		n6_idata_p0_30_ <= $random;
		n6_idata_p0_31_ <= $random;
		n6_idata_p0_32_ <= $random;
		n6_idata_p0_33_ <= $random;
		n6_idata_p0_34_ <= $random;
		n6_ivalid_p0 <= $random;
		n6_ivch_p0 <= $random;
		n7_idata_p0_0_ <= $random;
		n7_idata_p0_1_ <= $random;
		n7_idata_p0_2_ <= $random;
		n7_idata_p0_3_ <= $random;
		n7_idata_p0_4_ <= $random;
		n7_idata_p0_5_ <= $random;
		n7_idata_p0_6_ <= $random;
		n7_idata_p0_7_ <= $random;
		n7_idata_p0_8_ <= $random;
		n7_idata_p0_9_ <= $random;
		n7_idata_p0_10_ <= $random;
		n7_idata_p0_11_ <= $random;
		n7_idata_p0_12_ <= $random;
		n7_idata_p0_13_ <= $random;
		n7_idata_p0_14_ <= $random;
		n7_idata_p0_15_ <= $random;
		n7_idata_p0_16_ <= $random;
		n7_idata_p0_17_ <= $random;
		n7_idata_p0_18_ <= $random;
		n7_idata_p0_19_ <= $random;
		n7_idata_p0_20_ <= $random;
		n7_idata_p0_21_ <= $random;
		n7_idata_p0_22_ <= $random;
		n7_idata_p0_23_ <= $random;
		n7_idata_p0_24_ <= $random;
		n7_idata_p0_25_ <= $random;
		n7_idata_p0_26_ <= $random;
		n7_idata_p0_27_ <= $random;
		n7_idata_p0_28_ <= $random;
		n7_idata_p0_29_ <= $random;
		n7_idata_p0_30_ <= $random;
		n7_idata_p0_31_ <= $random;
		n7_idata_p0_32_ <= $random;
		n7_idata_p0_33_ <= $random;
		n7_idata_p0_34_ <= $random;
		n7_ivalid_p0 <= $random;
		n7_ivch_p0 <= $random;
		n8_idata_p0_0_ <= $random;
		n8_idata_p0_1_ <= $random;
		n8_idata_p0_2_ <= $random;
		n8_idata_p0_3_ <= $random;
		n8_idata_p0_4_ <= $random;
		n8_idata_p0_5_ <= $random;
		n8_idata_p0_6_ <= $random;
		n8_idata_p0_7_ <= $random;
		n8_idata_p0_8_ <= $random;
		n8_idata_p0_9_ <= $random;
		n8_idata_p0_10_ <= $random;
		n8_idata_p0_11_ <= $random;
		n8_idata_p0_12_ <= $random;
		n8_idata_p0_13_ <= $random;
		n8_idata_p0_14_ <= $random;
		n8_idata_p0_15_ <= $random;
		n8_idata_p0_16_ <= $random;
		n8_idata_p0_17_ <= $random;
		n8_idata_p0_18_ <= $random;
		n8_idata_p0_19_ <= $random;
		n8_idata_p0_20_ <= $random;
		n8_idata_p0_21_ <= $random;
		n8_idata_p0_22_ <= $random;
		n8_idata_p0_23_ <= $random;
		n8_idata_p0_24_ <= $random;
		n8_idata_p0_25_ <= $random;
		n8_idata_p0_26_ <= $random;
		n8_idata_p0_27_ <= $random;
		n8_idata_p0_28_ <= $random;
		n8_idata_p0_29_ <= $random;
		n8_idata_p0_30_ <= $random;
		n8_idata_p0_31_ <= $random;
		n8_idata_p0_32_ <= $random;
		n8_idata_p0_33_ <= $random;
		n8_idata_p0_34_ <= $random;
		n8_ivalid_p0 <= $random;
		n8_ivch_p0 <= $random;
		rst_ <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge clk[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else 
begin
			if(!(n0_ordy_p0_0__gfpga === n0_ordy_p0_0__bench) && !(n0_ordy_p0_0__bench === 1'bx)) begin
				n0_ordy_p0_0__flag <= 1'b1;
			end else begin
				n0_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n0_ordy_p0_1__gfpga === n0_ordy_p0_1__bench) && !(n0_ordy_p0_1__bench === 1'bx)) begin
				n0_ordy_p0_1__flag <= 1'b1;
			end else begin
				n0_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n0_odata_p0_0__gfpga === n0_odata_p0_0__bench) && !(n0_odata_p0_0__bench === 1'bx)) begin
				n0_odata_p0_0__flag <= 1'b1;
			end else begin
				n0_odata_p0_0__flag<= 1'b0;
			end
			if(!(n0_odata_p0_1__gfpga === n0_odata_p0_1__bench) && !(n0_odata_p0_1__bench === 1'bx)) begin
				n0_odata_p0_1__flag <= 1'b1;
			end else begin
				n0_odata_p0_1__flag<= 1'b0;
			end
			if(!(n0_odata_p0_2__gfpga === n0_odata_p0_2__bench) && !(n0_odata_p0_2__bench === 1'bx)) begin
				n0_odata_p0_2__flag <= 1'b1;
			end else begin
				n0_odata_p0_2__flag<= 1'b0;
			end
			if(!(n0_odata_p0_3__gfpga === n0_odata_p0_3__bench) && !(n0_odata_p0_3__bench === 1'bx)) begin
				n0_odata_p0_3__flag <= 1'b1;
			end else begin
				n0_odata_p0_3__flag<= 1'b0;
			end
			if(!(n0_odata_p0_4__gfpga === n0_odata_p0_4__bench) && !(n0_odata_p0_4__bench === 1'bx)) begin
				n0_odata_p0_4__flag <= 1'b1;
			end else begin
				n0_odata_p0_4__flag<= 1'b0;
			end
			if(!(n0_odata_p0_5__gfpga === n0_odata_p0_5__bench) && !(n0_odata_p0_5__bench === 1'bx)) begin
				n0_odata_p0_5__flag <= 1'b1;
			end else begin
				n0_odata_p0_5__flag<= 1'b0;
			end
			if(!(n0_odata_p0_6__gfpga === n0_odata_p0_6__bench) && !(n0_odata_p0_6__bench === 1'bx)) begin
				n0_odata_p0_6__flag <= 1'b1;
			end else begin
				n0_odata_p0_6__flag<= 1'b0;
			end
			if(!(n0_odata_p0_7__gfpga === n0_odata_p0_7__bench) && !(n0_odata_p0_7__bench === 1'bx)) begin
				n0_odata_p0_7__flag <= 1'b1;
			end else begin
				n0_odata_p0_7__flag<= 1'b0;
			end
			if(!(n0_odata_p0_8__gfpga === n0_odata_p0_8__bench) && !(n0_odata_p0_8__bench === 1'bx)) begin
				n0_odata_p0_8__flag <= 1'b1;
			end else begin
				n0_odata_p0_8__flag<= 1'b0;
			end
			if(!(n0_odata_p0_9__gfpga === n0_odata_p0_9__bench) && !(n0_odata_p0_9__bench === 1'bx)) begin
				n0_odata_p0_9__flag <= 1'b1;
			end else begin
				n0_odata_p0_9__flag<= 1'b0;
			end
			if(!(n0_odata_p0_10__gfpga === n0_odata_p0_10__bench) && !(n0_odata_p0_10__bench === 1'bx)) begin
				n0_odata_p0_10__flag <= 1'b1;
			end else begin
				n0_odata_p0_10__flag<= 1'b0;
			end
			if(!(n0_odata_p0_11__gfpga === n0_odata_p0_11__bench) && !(n0_odata_p0_11__bench === 1'bx)) begin
				n0_odata_p0_11__flag <= 1'b1;
			end else begin
				n0_odata_p0_11__flag<= 1'b0;
			end
			if(!(n0_odata_p0_12__gfpga === n0_odata_p0_12__bench) && !(n0_odata_p0_12__bench === 1'bx)) begin
				n0_odata_p0_12__flag <= 1'b1;
			end else begin
				n0_odata_p0_12__flag<= 1'b0;
			end
			if(!(n0_odata_p0_13__gfpga === n0_odata_p0_13__bench) && !(n0_odata_p0_13__bench === 1'bx)) begin
				n0_odata_p0_13__flag <= 1'b1;
			end else begin
				n0_odata_p0_13__flag<= 1'b0;
			end
			if(!(n0_odata_p0_14__gfpga === n0_odata_p0_14__bench) && !(n0_odata_p0_14__bench === 1'bx)) begin
				n0_odata_p0_14__flag <= 1'b1;
			end else begin
				n0_odata_p0_14__flag<= 1'b0;
			end
			if(!(n0_odata_p0_15__gfpga === n0_odata_p0_15__bench) && !(n0_odata_p0_15__bench === 1'bx)) begin
				n0_odata_p0_15__flag <= 1'b1;
			end else begin
				n0_odata_p0_15__flag<= 1'b0;
			end
			if(!(n0_odata_p0_16__gfpga === n0_odata_p0_16__bench) && !(n0_odata_p0_16__bench === 1'bx)) begin
				n0_odata_p0_16__flag <= 1'b1;
			end else begin
				n0_odata_p0_16__flag<= 1'b0;
			end
			if(!(n0_odata_p0_17__gfpga === n0_odata_p0_17__bench) && !(n0_odata_p0_17__bench === 1'bx)) begin
				n0_odata_p0_17__flag <= 1'b1;
			end else begin
				n0_odata_p0_17__flag<= 1'b0;
			end
			if(!(n0_odata_p0_18__gfpga === n0_odata_p0_18__bench) && !(n0_odata_p0_18__bench === 1'bx)) begin
				n0_odata_p0_18__flag <= 1'b1;
			end else begin
				n0_odata_p0_18__flag<= 1'b0;
			end
			if(!(n0_odata_p0_19__gfpga === n0_odata_p0_19__bench) && !(n0_odata_p0_19__bench === 1'bx)) begin
				n0_odata_p0_19__flag <= 1'b1;
			end else begin
				n0_odata_p0_19__flag<= 1'b0;
			end
			if(!(n0_odata_p0_20__gfpga === n0_odata_p0_20__bench) && !(n0_odata_p0_20__bench === 1'bx)) begin
				n0_odata_p0_20__flag <= 1'b1;
			end else begin
				n0_odata_p0_20__flag<= 1'b0;
			end
			if(!(n0_odata_p0_21__gfpga === n0_odata_p0_21__bench) && !(n0_odata_p0_21__bench === 1'bx)) begin
				n0_odata_p0_21__flag <= 1'b1;
			end else begin
				n0_odata_p0_21__flag<= 1'b0;
			end
			if(!(n0_odata_p0_22__gfpga === n0_odata_p0_22__bench) && !(n0_odata_p0_22__bench === 1'bx)) begin
				n0_odata_p0_22__flag <= 1'b1;
			end else begin
				n0_odata_p0_22__flag<= 1'b0;
			end
			if(!(n0_odata_p0_23__gfpga === n0_odata_p0_23__bench) && !(n0_odata_p0_23__bench === 1'bx)) begin
				n0_odata_p0_23__flag <= 1'b1;
			end else begin
				n0_odata_p0_23__flag<= 1'b0;
			end
			if(!(n0_odata_p0_24__gfpga === n0_odata_p0_24__bench) && !(n0_odata_p0_24__bench === 1'bx)) begin
				n0_odata_p0_24__flag <= 1'b1;
			end else begin
				n0_odata_p0_24__flag<= 1'b0;
			end
			if(!(n0_odata_p0_25__gfpga === n0_odata_p0_25__bench) && !(n0_odata_p0_25__bench === 1'bx)) begin
				n0_odata_p0_25__flag <= 1'b1;
			end else begin
				n0_odata_p0_25__flag<= 1'b0;
			end
			if(!(n0_odata_p0_26__gfpga === n0_odata_p0_26__bench) && !(n0_odata_p0_26__bench === 1'bx)) begin
				n0_odata_p0_26__flag <= 1'b1;
			end else begin
				n0_odata_p0_26__flag<= 1'b0;
			end
			if(!(n0_odata_p0_27__gfpga === n0_odata_p0_27__bench) && !(n0_odata_p0_27__bench === 1'bx)) begin
				n0_odata_p0_27__flag <= 1'b1;
			end else begin
				n0_odata_p0_27__flag<= 1'b0;
			end
			if(!(n0_odata_p0_28__gfpga === n0_odata_p0_28__bench) && !(n0_odata_p0_28__bench === 1'bx)) begin
				n0_odata_p0_28__flag <= 1'b1;
			end else begin
				n0_odata_p0_28__flag<= 1'b0;
			end
			if(!(n0_odata_p0_29__gfpga === n0_odata_p0_29__bench) && !(n0_odata_p0_29__bench === 1'bx)) begin
				n0_odata_p0_29__flag <= 1'b1;
			end else begin
				n0_odata_p0_29__flag<= 1'b0;
			end
			if(!(n0_odata_p0_30__gfpga === n0_odata_p0_30__bench) && !(n0_odata_p0_30__bench === 1'bx)) begin
				n0_odata_p0_30__flag <= 1'b1;
			end else begin
				n0_odata_p0_30__flag<= 1'b0;
			end
			if(!(n0_odata_p0_31__gfpga === n0_odata_p0_31__bench) && !(n0_odata_p0_31__bench === 1'bx)) begin
				n0_odata_p0_31__flag <= 1'b1;
			end else begin
				n0_odata_p0_31__flag<= 1'b0;
			end
			if(!(n0_odata_p0_32__gfpga === n0_odata_p0_32__bench) && !(n0_odata_p0_32__bench === 1'bx)) begin
				n0_odata_p0_32__flag <= 1'b1;
			end else begin
				n0_odata_p0_32__flag<= 1'b0;
			end
			if(!(n0_odata_p0_33__gfpga === n0_odata_p0_33__bench) && !(n0_odata_p0_33__bench === 1'bx)) begin
				n0_odata_p0_33__flag <= 1'b1;
			end else begin
				n0_odata_p0_33__flag<= 1'b0;
			end
			if(!(n0_odata_p0_34__gfpga === n0_odata_p0_34__bench) && !(n0_odata_p0_34__bench === 1'bx)) begin
				n0_odata_p0_34__flag <= 1'b1;
			end else begin
				n0_odata_p0_34__flag<= 1'b0;
			end
			if(!(n0_ovalid_p0_gfpga === n0_ovalid_p0_bench) && !(n0_ovalid_p0_bench === 1'bx)) begin
				n0_ovalid_p0_flag <= 1'b1;
			end else begin
				n0_ovalid_p0_flag<= 1'b0;
			end
			if(!(n1_ordy_p0_0__gfpga === n1_ordy_p0_0__bench) && !(n1_ordy_p0_0__bench === 1'bx)) begin
				n1_ordy_p0_0__flag <= 1'b1;
			end else begin
				n1_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n1_ordy_p0_1__gfpga === n1_ordy_p0_1__bench) && !(n1_ordy_p0_1__bench === 1'bx)) begin
				n1_ordy_p0_1__flag <= 1'b1;
			end else begin
				n1_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n1_odata_p0_0__gfpga === n1_odata_p0_0__bench) && !(n1_odata_p0_0__bench === 1'bx)) begin
				n1_odata_p0_0__flag <= 1'b1;
			end else begin
				n1_odata_p0_0__flag<= 1'b0;
			end
			if(!(n1_odata_p0_1__gfpga === n1_odata_p0_1__bench) && !(n1_odata_p0_1__bench === 1'bx)) begin
				n1_odata_p0_1__flag <= 1'b1;
			end else begin
				n1_odata_p0_1__flag<= 1'b0;
			end
			if(!(n1_odata_p0_2__gfpga === n1_odata_p0_2__bench) && !(n1_odata_p0_2__bench === 1'bx)) begin
				n1_odata_p0_2__flag <= 1'b1;
			end else begin
				n1_odata_p0_2__flag<= 1'b0;
			end
			if(!(n1_odata_p0_3__gfpga === n1_odata_p0_3__bench) && !(n1_odata_p0_3__bench === 1'bx)) begin
				n1_odata_p0_3__flag <= 1'b1;
			end else begin
				n1_odata_p0_3__flag<= 1'b0;
			end
			if(!(n1_odata_p0_4__gfpga === n1_odata_p0_4__bench) && !(n1_odata_p0_4__bench === 1'bx)) begin
				n1_odata_p0_4__flag <= 1'b1;
			end else begin
				n1_odata_p0_4__flag<= 1'b0;
			end
			if(!(n1_odata_p0_5__gfpga === n1_odata_p0_5__bench) && !(n1_odata_p0_5__bench === 1'bx)) begin
				n1_odata_p0_5__flag <= 1'b1;
			end else begin
				n1_odata_p0_5__flag<= 1'b0;
			end
			if(!(n1_odata_p0_6__gfpga === n1_odata_p0_6__bench) && !(n1_odata_p0_6__bench === 1'bx)) begin
				n1_odata_p0_6__flag <= 1'b1;
			end else begin
				n1_odata_p0_6__flag<= 1'b0;
			end
			if(!(n1_odata_p0_7__gfpga === n1_odata_p0_7__bench) && !(n1_odata_p0_7__bench === 1'bx)) begin
				n1_odata_p0_7__flag <= 1'b1;
			end else begin
				n1_odata_p0_7__flag<= 1'b0;
			end
			if(!(n1_odata_p0_8__gfpga === n1_odata_p0_8__bench) && !(n1_odata_p0_8__bench === 1'bx)) begin
				n1_odata_p0_8__flag <= 1'b1;
			end else begin
				n1_odata_p0_8__flag<= 1'b0;
			end
			if(!(n1_odata_p0_9__gfpga === n1_odata_p0_9__bench) && !(n1_odata_p0_9__bench === 1'bx)) begin
				n1_odata_p0_9__flag <= 1'b1;
			end else begin
				n1_odata_p0_9__flag<= 1'b0;
			end
			if(!(n1_odata_p0_10__gfpga === n1_odata_p0_10__bench) && !(n1_odata_p0_10__bench === 1'bx)) begin
				n1_odata_p0_10__flag <= 1'b1;
			end else begin
				n1_odata_p0_10__flag<= 1'b0;
			end
			if(!(n1_odata_p0_11__gfpga === n1_odata_p0_11__bench) && !(n1_odata_p0_11__bench === 1'bx)) begin
				n1_odata_p0_11__flag <= 1'b1;
			end else begin
				n1_odata_p0_11__flag<= 1'b0;
			end
			if(!(n1_odata_p0_12__gfpga === n1_odata_p0_12__bench) && !(n1_odata_p0_12__bench === 1'bx)) begin
				n1_odata_p0_12__flag <= 1'b1;
			end else begin
				n1_odata_p0_12__flag<= 1'b0;
			end
			if(!(n1_odata_p0_13__gfpga === n1_odata_p0_13__bench) && !(n1_odata_p0_13__bench === 1'bx)) begin
				n1_odata_p0_13__flag <= 1'b1;
			end else begin
				n1_odata_p0_13__flag<= 1'b0;
			end
			if(!(n1_odata_p0_14__gfpga === n1_odata_p0_14__bench) && !(n1_odata_p0_14__bench === 1'bx)) begin
				n1_odata_p0_14__flag <= 1'b1;
			end else begin
				n1_odata_p0_14__flag<= 1'b0;
			end
			if(!(n1_odata_p0_15__gfpga === n1_odata_p0_15__bench) && !(n1_odata_p0_15__bench === 1'bx)) begin
				n1_odata_p0_15__flag <= 1'b1;
			end else begin
				n1_odata_p0_15__flag<= 1'b0;
			end
			if(!(n1_odata_p0_16__gfpga === n1_odata_p0_16__bench) && !(n1_odata_p0_16__bench === 1'bx)) begin
				n1_odata_p0_16__flag <= 1'b1;
			end else begin
				n1_odata_p0_16__flag<= 1'b0;
			end
			if(!(n1_odata_p0_17__gfpga === n1_odata_p0_17__bench) && !(n1_odata_p0_17__bench === 1'bx)) begin
				n1_odata_p0_17__flag <= 1'b1;
			end else begin
				n1_odata_p0_17__flag<= 1'b0;
			end
			if(!(n1_odata_p0_18__gfpga === n1_odata_p0_18__bench) && !(n1_odata_p0_18__bench === 1'bx)) begin
				n1_odata_p0_18__flag <= 1'b1;
			end else begin
				n1_odata_p0_18__flag<= 1'b0;
			end
			if(!(n1_odata_p0_19__gfpga === n1_odata_p0_19__bench) && !(n1_odata_p0_19__bench === 1'bx)) begin
				n1_odata_p0_19__flag <= 1'b1;
			end else begin
				n1_odata_p0_19__flag<= 1'b0;
			end
			if(!(n1_odata_p0_20__gfpga === n1_odata_p0_20__bench) && !(n1_odata_p0_20__bench === 1'bx)) begin
				n1_odata_p0_20__flag <= 1'b1;
			end else begin
				n1_odata_p0_20__flag<= 1'b0;
			end
			if(!(n1_odata_p0_21__gfpga === n1_odata_p0_21__bench) && !(n1_odata_p0_21__bench === 1'bx)) begin
				n1_odata_p0_21__flag <= 1'b1;
			end else begin
				n1_odata_p0_21__flag<= 1'b0;
			end
			if(!(n1_odata_p0_22__gfpga === n1_odata_p0_22__bench) && !(n1_odata_p0_22__bench === 1'bx)) begin
				n1_odata_p0_22__flag <= 1'b1;
			end else begin
				n1_odata_p0_22__flag<= 1'b0;
			end
			if(!(n1_odata_p0_23__gfpga === n1_odata_p0_23__bench) && !(n1_odata_p0_23__bench === 1'bx)) begin
				n1_odata_p0_23__flag <= 1'b1;
			end else begin
				n1_odata_p0_23__flag<= 1'b0;
			end
			if(!(n1_odata_p0_24__gfpga === n1_odata_p0_24__bench) && !(n1_odata_p0_24__bench === 1'bx)) begin
				n1_odata_p0_24__flag <= 1'b1;
			end else begin
				n1_odata_p0_24__flag<= 1'b0;
			end
			if(!(n1_odata_p0_25__gfpga === n1_odata_p0_25__bench) && !(n1_odata_p0_25__bench === 1'bx)) begin
				n1_odata_p0_25__flag <= 1'b1;
			end else begin
				n1_odata_p0_25__flag<= 1'b0;
			end
			if(!(n1_odata_p0_26__gfpga === n1_odata_p0_26__bench) && !(n1_odata_p0_26__bench === 1'bx)) begin
				n1_odata_p0_26__flag <= 1'b1;
			end else begin
				n1_odata_p0_26__flag<= 1'b0;
			end
			if(!(n1_odata_p0_27__gfpga === n1_odata_p0_27__bench) && !(n1_odata_p0_27__bench === 1'bx)) begin
				n1_odata_p0_27__flag <= 1'b1;
			end else begin
				n1_odata_p0_27__flag<= 1'b0;
			end
			if(!(n1_odata_p0_28__gfpga === n1_odata_p0_28__bench) && !(n1_odata_p0_28__bench === 1'bx)) begin
				n1_odata_p0_28__flag <= 1'b1;
			end else begin
				n1_odata_p0_28__flag<= 1'b0;
			end
			if(!(n1_odata_p0_29__gfpga === n1_odata_p0_29__bench) && !(n1_odata_p0_29__bench === 1'bx)) begin
				n1_odata_p0_29__flag <= 1'b1;
			end else begin
				n1_odata_p0_29__flag<= 1'b0;
			end
			if(!(n1_odata_p0_30__gfpga === n1_odata_p0_30__bench) && !(n1_odata_p0_30__bench === 1'bx)) begin
				n1_odata_p0_30__flag <= 1'b1;
			end else begin
				n1_odata_p0_30__flag<= 1'b0;
			end
			if(!(n1_odata_p0_31__gfpga === n1_odata_p0_31__bench) && !(n1_odata_p0_31__bench === 1'bx)) begin
				n1_odata_p0_31__flag <= 1'b1;
			end else begin
				n1_odata_p0_31__flag<= 1'b0;
			end
			if(!(n1_odata_p0_32__gfpga === n1_odata_p0_32__bench) && !(n1_odata_p0_32__bench === 1'bx)) begin
				n1_odata_p0_32__flag <= 1'b1;
			end else begin
				n1_odata_p0_32__flag<= 1'b0;
			end
			if(!(n1_odata_p0_33__gfpga === n1_odata_p0_33__bench) && !(n1_odata_p0_33__bench === 1'bx)) begin
				n1_odata_p0_33__flag <= 1'b1;
			end else begin
				n1_odata_p0_33__flag<= 1'b0;
			end
			if(!(n1_odata_p0_34__gfpga === n1_odata_p0_34__bench) && !(n1_odata_p0_34__bench === 1'bx)) begin
				n1_odata_p0_34__flag <= 1'b1;
			end else begin
				n1_odata_p0_34__flag<= 1'b0;
			end
			if(!(n1_ovalid_p0_gfpga === n1_ovalid_p0_bench) && !(n1_ovalid_p0_bench === 1'bx)) begin
				n1_ovalid_p0_flag <= 1'b1;
			end else begin
				n1_ovalid_p0_flag<= 1'b0;
			end
			if(!(n2_ordy_p0_0__gfpga === n2_ordy_p0_0__bench) && !(n2_ordy_p0_0__bench === 1'bx)) begin
				n2_ordy_p0_0__flag <= 1'b1;
			end else begin
				n2_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n2_ordy_p0_1__gfpga === n2_ordy_p0_1__bench) && !(n2_ordy_p0_1__bench === 1'bx)) begin
				n2_ordy_p0_1__flag <= 1'b1;
			end else begin
				n2_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n2_odata_p0_0__gfpga === n2_odata_p0_0__bench) && !(n2_odata_p0_0__bench === 1'bx)) begin
				n2_odata_p0_0__flag <= 1'b1;
			end else begin
				n2_odata_p0_0__flag<= 1'b0;
			end
			if(!(n2_odata_p0_1__gfpga === n2_odata_p0_1__bench) && !(n2_odata_p0_1__bench === 1'bx)) begin
				n2_odata_p0_1__flag <= 1'b1;
			end else begin
				n2_odata_p0_1__flag<= 1'b0;
			end
			if(!(n2_odata_p0_2__gfpga === n2_odata_p0_2__bench) && !(n2_odata_p0_2__bench === 1'bx)) begin
				n2_odata_p0_2__flag <= 1'b1;
			end else begin
				n2_odata_p0_2__flag<= 1'b0;
			end
			if(!(n2_odata_p0_3__gfpga === n2_odata_p0_3__bench) && !(n2_odata_p0_3__bench === 1'bx)) begin
				n2_odata_p0_3__flag <= 1'b1;
			end else begin
				n2_odata_p0_3__flag<= 1'b0;
			end
			if(!(n2_odata_p0_4__gfpga === n2_odata_p0_4__bench) && !(n2_odata_p0_4__bench === 1'bx)) begin
				n2_odata_p0_4__flag <= 1'b1;
			end else begin
				n2_odata_p0_4__flag<= 1'b0;
			end
			if(!(n2_odata_p0_5__gfpga === n2_odata_p0_5__bench) && !(n2_odata_p0_5__bench === 1'bx)) begin
				n2_odata_p0_5__flag <= 1'b1;
			end else begin
				n2_odata_p0_5__flag<= 1'b0;
			end
			if(!(n2_odata_p0_6__gfpga === n2_odata_p0_6__bench) && !(n2_odata_p0_6__bench === 1'bx)) begin
				n2_odata_p0_6__flag <= 1'b1;
			end else begin
				n2_odata_p0_6__flag<= 1'b0;
			end
			if(!(n2_odata_p0_7__gfpga === n2_odata_p0_7__bench) && !(n2_odata_p0_7__bench === 1'bx)) begin
				n2_odata_p0_7__flag <= 1'b1;
			end else begin
				n2_odata_p0_7__flag<= 1'b0;
			end
			if(!(n2_odata_p0_8__gfpga === n2_odata_p0_8__bench) && !(n2_odata_p0_8__bench === 1'bx)) begin
				n2_odata_p0_8__flag <= 1'b1;
			end else begin
				n2_odata_p0_8__flag<= 1'b0;
			end
			if(!(n2_odata_p0_9__gfpga === n2_odata_p0_9__bench) && !(n2_odata_p0_9__bench === 1'bx)) begin
				n2_odata_p0_9__flag <= 1'b1;
			end else begin
				n2_odata_p0_9__flag<= 1'b0;
			end
			if(!(n2_odata_p0_10__gfpga === n2_odata_p0_10__bench) && !(n2_odata_p0_10__bench === 1'bx)) begin
				n2_odata_p0_10__flag <= 1'b1;
			end else begin
				n2_odata_p0_10__flag<= 1'b0;
			end
			if(!(n2_odata_p0_11__gfpga === n2_odata_p0_11__bench) && !(n2_odata_p0_11__bench === 1'bx)) begin
				n2_odata_p0_11__flag <= 1'b1;
			end else begin
				n2_odata_p0_11__flag<= 1'b0;
			end
			if(!(n2_odata_p0_12__gfpga === n2_odata_p0_12__bench) && !(n2_odata_p0_12__bench === 1'bx)) begin
				n2_odata_p0_12__flag <= 1'b1;
			end else begin
				n2_odata_p0_12__flag<= 1'b0;
			end
			if(!(n2_odata_p0_13__gfpga === n2_odata_p0_13__bench) && !(n2_odata_p0_13__bench === 1'bx)) begin
				n2_odata_p0_13__flag <= 1'b1;
			end else begin
				n2_odata_p0_13__flag<= 1'b0;
			end
			if(!(n2_odata_p0_14__gfpga === n2_odata_p0_14__bench) && !(n2_odata_p0_14__bench === 1'bx)) begin
				n2_odata_p0_14__flag <= 1'b1;
			end else begin
				n2_odata_p0_14__flag<= 1'b0;
			end
			if(!(n2_odata_p0_15__gfpga === n2_odata_p0_15__bench) && !(n2_odata_p0_15__bench === 1'bx)) begin
				n2_odata_p0_15__flag <= 1'b1;
			end else begin
				n2_odata_p0_15__flag<= 1'b0;
			end
			if(!(n2_odata_p0_16__gfpga === n2_odata_p0_16__bench) && !(n2_odata_p0_16__bench === 1'bx)) begin
				n2_odata_p0_16__flag <= 1'b1;
			end else begin
				n2_odata_p0_16__flag<= 1'b0;
			end
			if(!(n2_odata_p0_17__gfpga === n2_odata_p0_17__bench) && !(n2_odata_p0_17__bench === 1'bx)) begin
				n2_odata_p0_17__flag <= 1'b1;
			end else begin
				n2_odata_p0_17__flag<= 1'b0;
			end
			if(!(n2_odata_p0_18__gfpga === n2_odata_p0_18__bench) && !(n2_odata_p0_18__bench === 1'bx)) begin
				n2_odata_p0_18__flag <= 1'b1;
			end else begin
				n2_odata_p0_18__flag<= 1'b0;
			end
			if(!(n2_odata_p0_19__gfpga === n2_odata_p0_19__bench) && !(n2_odata_p0_19__bench === 1'bx)) begin
				n2_odata_p0_19__flag <= 1'b1;
			end else begin
				n2_odata_p0_19__flag<= 1'b0;
			end
			if(!(n2_odata_p0_20__gfpga === n2_odata_p0_20__bench) && !(n2_odata_p0_20__bench === 1'bx)) begin
				n2_odata_p0_20__flag <= 1'b1;
			end else begin
				n2_odata_p0_20__flag<= 1'b0;
			end
			if(!(n2_odata_p0_21__gfpga === n2_odata_p0_21__bench) && !(n2_odata_p0_21__bench === 1'bx)) begin
				n2_odata_p0_21__flag <= 1'b1;
			end else begin
				n2_odata_p0_21__flag<= 1'b0;
			end
			if(!(n2_odata_p0_22__gfpga === n2_odata_p0_22__bench) && !(n2_odata_p0_22__bench === 1'bx)) begin
				n2_odata_p0_22__flag <= 1'b1;
			end else begin
				n2_odata_p0_22__flag<= 1'b0;
			end
			if(!(n2_odata_p0_23__gfpga === n2_odata_p0_23__bench) && !(n2_odata_p0_23__bench === 1'bx)) begin
				n2_odata_p0_23__flag <= 1'b1;
			end else begin
				n2_odata_p0_23__flag<= 1'b0;
			end
			if(!(n2_odata_p0_24__gfpga === n2_odata_p0_24__bench) && !(n2_odata_p0_24__bench === 1'bx)) begin
				n2_odata_p0_24__flag <= 1'b1;
			end else begin
				n2_odata_p0_24__flag<= 1'b0;
			end
			if(!(n2_odata_p0_25__gfpga === n2_odata_p0_25__bench) && !(n2_odata_p0_25__bench === 1'bx)) begin
				n2_odata_p0_25__flag <= 1'b1;
			end else begin
				n2_odata_p0_25__flag<= 1'b0;
			end
			if(!(n2_odata_p0_26__gfpga === n2_odata_p0_26__bench) && !(n2_odata_p0_26__bench === 1'bx)) begin
				n2_odata_p0_26__flag <= 1'b1;
			end else begin
				n2_odata_p0_26__flag<= 1'b0;
			end
			if(!(n2_odata_p0_27__gfpga === n2_odata_p0_27__bench) && !(n2_odata_p0_27__bench === 1'bx)) begin
				n2_odata_p0_27__flag <= 1'b1;
			end else begin
				n2_odata_p0_27__flag<= 1'b0;
			end
			if(!(n2_odata_p0_28__gfpga === n2_odata_p0_28__bench) && !(n2_odata_p0_28__bench === 1'bx)) begin
				n2_odata_p0_28__flag <= 1'b1;
			end else begin
				n2_odata_p0_28__flag<= 1'b0;
			end
			if(!(n2_odata_p0_29__gfpga === n2_odata_p0_29__bench) && !(n2_odata_p0_29__bench === 1'bx)) begin
				n2_odata_p0_29__flag <= 1'b1;
			end else begin
				n2_odata_p0_29__flag<= 1'b0;
			end
			if(!(n2_odata_p0_30__gfpga === n2_odata_p0_30__bench) && !(n2_odata_p0_30__bench === 1'bx)) begin
				n2_odata_p0_30__flag <= 1'b1;
			end else begin
				n2_odata_p0_30__flag<= 1'b0;
			end
			if(!(n2_odata_p0_31__gfpga === n2_odata_p0_31__bench) && !(n2_odata_p0_31__bench === 1'bx)) begin
				n2_odata_p0_31__flag <= 1'b1;
			end else begin
				n2_odata_p0_31__flag<= 1'b0;
			end
			if(!(n2_odata_p0_32__gfpga === n2_odata_p0_32__bench) && !(n2_odata_p0_32__bench === 1'bx)) begin
				n2_odata_p0_32__flag <= 1'b1;
			end else begin
				n2_odata_p0_32__flag<= 1'b0;
			end
			if(!(n2_odata_p0_33__gfpga === n2_odata_p0_33__bench) && !(n2_odata_p0_33__bench === 1'bx)) begin
				n2_odata_p0_33__flag <= 1'b1;
			end else begin
				n2_odata_p0_33__flag<= 1'b0;
			end
			if(!(n2_odata_p0_34__gfpga === n2_odata_p0_34__bench) && !(n2_odata_p0_34__bench === 1'bx)) begin
				n2_odata_p0_34__flag <= 1'b1;
			end else begin
				n2_odata_p0_34__flag<= 1'b0;
			end
			if(!(n2_ovalid_p0_gfpga === n2_ovalid_p0_bench) && !(n2_ovalid_p0_bench === 1'bx)) begin
				n2_ovalid_p0_flag <= 1'b1;
			end else begin
				n2_ovalid_p0_flag<= 1'b0;
			end
			if(!(n3_ordy_p0_0__gfpga === n3_ordy_p0_0__bench) && !(n3_ordy_p0_0__bench === 1'bx)) begin
				n3_ordy_p0_0__flag <= 1'b1;
			end else begin
				n3_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n3_ordy_p0_1__gfpga === n3_ordy_p0_1__bench) && !(n3_ordy_p0_1__bench === 1'bx)) begin
				n3_ordy_p0_1__flag <= 1'b1;
			end else begin
				n3_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n3_odata_p0_0__gfpga === n3_odata_p0_0__bench) && !(n3_odata_p0_0__bench === 1'bx)) begin
				n3_odata_p0_0__flag <= 1'b1;
			end else begin
				n3_odata_p0_0__flag<= 1'b0;
			end
			if(!(n3_odata_p0_1__gfpga === n3_odata_p0_1__bench) && !(n3_odata_p0_1__bench === 1'bx)) begin
				n3_odata_p0_1__flag <= 1'b1;
			end else begin
				n3_odata_p0_1__flag<= 1'b0;
			end
			if(!(n3_odata_p0_2__gfpga === n3_odata_p0_2__bench) && !(n3_odata_p0_2__bench === 1'bx)) begin
				n3_odata_p0_2__flag <= 1'b1;
			end else begin
				n3_odata_p0_2__flag<= 1'b0;
			end
			if(!(n3_odata_p0_3__gfpga === n3_odata_p0_3__bench) && !(n3_odata_p0_3__bench === 1'bx)) begin
				n3_odata_p0_3__flag <= 1'b1;
			end else begin
				n3_odata_p0_3__flag<= 1'b0;
			end
			if(!(n3_odata_p0_4__gfpga === n3_odata_p0_4__bench) && !(n3_odata_p0_4__bench === 1'bx)) begin
				n3_odata_p0_4__flag <= 1'b1;
			end else begin
				n3_odata_p0_4__flag<= 1'b0;
			end
			if(!(n3_odata_p0_5__gfpga === n3_odata_p0_5__bench) && !(n3_odata_p0_5__bench === 1'bx)) begin
				n3_odata_p0_5__flag <= 1'b1;
			end else begin
				n3_odata_p0_5__flag<= 1'b0;
			end
			if(!(n3_odata_p0_6__gfpga === n3_odata_p0_6__bench) && !(n3_odata_p0_6__bench === 1'bx)) begin
				n3_odata_p0_6__flag <= 1'b1;
			end else begin
				n3_odata_p0_6__flag<= 1'b0;
			end
			if(!(n3_odata_p0_7__gfpga === n3_odata_p0_7__bench) && !(n3_odata_p0_7__bench === 1'bx)) begin
				n3_odata_p0_7__flag <= 1'b1;
			end else begin
				n3_odata_p0_7__flag<= 1'b0;
			end
			if(!(n3_odata_p0_8__gfpga === n3_odata_p0_8__bench) && !(n3_odata_p0_8__bench === 1'bx)) begin
				n3_odata_p0_8__flag <= 1'b1;
			end else begin
				n3_odata_p0_8__flag<= 1'b0;
			end
			if(!(n3_odata_p0_9__gfpga === n3_odata_p0_9__bench) && !(n3_odata_p0_9__bench === 1'bx)) begin
				n3_odata_p0_9__flag <= 1'b1;
			end else begin
				n3_odata_p0_9__flag<= 1'b0;
			end
			if(!(n3_odata_p0_10__gfpga === n3_odata_p0_10__bench) && !(n3_odata_p0_10__bench === 1'bx)) begin
				n3_odata_p0_10__flag <= 1'b1;
			end else begin
				n3_odata_p0_10__flag<= 1'b0;
			end
			if(!(n3_odata_p0_11__gfpga === n3_odata_p0_11__bench) && !(n3_odata_p0_11__bench === 1'bx)) begin
				n3_odata_p0_11__flag <= 1'b1;
			end else begin
				n3_odata_p0_11__flag<= 1'b0;
			end
			if(!(n3_odata_p0_12__gfpga === n3_odata_p0_12__bench) && !(n3_odata_p0_12__bench === 1'bx)) begin
				n3_odata_p0_12__flag <= 1'b1;
			end else begin
				n3_odata_p0_12__flag<= 1'b0;
			end
			if(!(n3_odata_p0_13__gfpga === n3_odata_p0_13__bench) && !(n3_odata_p0_13__bench === 1'bx)) begin
				n3_odata_p0_13__flag <= 1'b1;
			end else begin
				n3_odata_p0_13__flag<= 1'b0;
			end
			if(!(n3_odata_p0_14__gfpga === n3_odata_p0_14__bench) && !(n3_odata_p0_14__bench === 1'bx)) begin
				n3_odata_p0_14__flag <= 1'b1;
			end else begin
				n3_odata_p0_14__flag<= 1'b0;
			end
			if(!(n3_odata_p0_15__gfpga === n3_odata_p0_15__bench) && !(n3_odata_p0_15__bench === 1'bx)) begin
				n3_odata_p0_15__flag <= 1'b1;
			end else begin
				n3_odata_p0_15__flag<= 1'b0;
			end
			if(!(n3_odata_p0_16__gfpga === n3_odata_p0_16__bench) && !(n3_odata_p0_16__bench === 1'bx)) begin
				n3_odata_p0_16__flag <= 1'b1;
			end else begin
				n3_odata_p0_16__flag<= 1'b0;
			end
			if(!(n3_odata_p0_17__gfpga === n3_odata_p0_17__bench) && !(n3_odata_p0_17__bench === 1'bx)) begin
				n3_odata_p0_17__flag <= 1'b1;
			end else begin
				n3_odata_p0_17__flag<= 1'b0;
			end
			if(!(n3_odata_p0_18__gfpga === n3_odata_p0_18__bench) && !(n3_odata_p0_18__bench === 1'bx)) begin
				n3_odata_p0_18__flag <= 1'b1;
			end else begin
				n3_odata_p0_18__flag<= 1'b0;
			end
			if(!(n3_odata_p0_19__gfpga === n3_odata_p0_19__bench) && !(n3_odata_p0_19__bench === 1'bx)) begin
				n3_odata_p0_19__flag <= 1'b1;
			end else begin
				n3_odata_p0_19__flag<= 1'b0;
			end
			if(!(n3_odata_p0_20__gfpga === n3_odata_p0_20__bench) && !(n3_odata_p0_20__bench === 1'bx)) begin
				n3_odata_p0_20__flag <= 1'b1;
			end else begin
				n3_odata_p0_20__flag<= 1'b0;
			end
			if(!(n3_odata_p0_21__gfpga === n3_odata_p0_21__bench) && !(n3_odata_p0_21__bench === 1'bx)) begin
				n3_odata_p0_21__flag <= 1'b1;
			end else begin
				n3_odata_p0_21__flag<= 1'b0;
			end
			if(!(n3_odata_p0_22__gfpga === n3_odata_p0_22__bench) && !(n3_odata_p0_22__bench === 1'bx)) begin
				n3_odata_p0_22__flag <= 1'b1;
			end else begin
				n3_odata_p0_22__flag<= 1'b0;
			end
			if(!(n3_odata_p0_23__gfpga === n3_odata_p0_23__bench) && !(n3_odata_p0_23__bench === 1'bx)) begin
				n3_odata_p0_23__flag <= 1'b1;
			end else begin
				n3_odata_p0_23__flag<= 1'b0;
			end
			if(!(n3_odata_p0_24__gfpga === n3_odata_p0_24__bench) && !(n3_odata_p0_24__bench === 1'bx)) begin
				n3_odata_p0_24__flag <= 1'b1;
			end else begin
				n3_odata_p0_24__flag<= 1'b0;
			end
			if(!(n3_odata_p0_25__gfpga === n3_odata_p0_25__bench) && !(n3_odata_p0_25__bench === 1'bx)) begin
				n3_odata_p0_25__flag <= 1'b1;
			end else begin
				n3_odata_p0_25__flag<= 1'b0;
			end
			if(!(n3_odata_p0_26__gfpga === n3_odata_p0_26__bench) && !(n3_odata_p0_26__bench === 1'bx)) begin
				n3_odata_p0_26__flag <= 1'b1;
			end else begin
				n3_odata_p0_26__flag<= 1'b0;
			end
			if(!(n3_odata_p0_27__gfpga === n3_odata_p0_27__bench) && !(n3_odata_p0_27__bench === 1'bx)) begin
				n3_odata_p0_27__flag <= 1'b1;
			end else begin
				n3_odata_p0_27__flag<= 1'b0;
			end
			if(!(n3_odata_p0_28__gfpga === n3_odata_p0_28__bench) && !(n3_odata_p0_28__bench === 1'bx)) begin
				n3_odata_p0_28__flag <= 1'b1;
			end else begin
				n3_odata_p0_28__flag<= 1'b0;
			end
			if(!(n3_odata_p0_29__gfpga === n3_odata_p0_29__bench) && !(n3_odata_p0_29__bench === 1'bx)) begin
				n3_odata_p0_29__flag <= 1'b1;
			end else begin
				n3_odata_p0_29__flag<= 1'b0;
			end
			if(!(n3_odata_p0_30__gfpga === n3_odata_p0_30__bench) && !(n3_odata_p0_30__bench === 1'bx)) begin
				n3_odata_p0_30__flag <= 1'b1;
			end else begin
				n3_odata_p0_30__flag<= 1'b0;
			end
			if(!(n3_odata_p0_31__gfpga === n3_odata_p0_31__bench) && !(n3_odata_p0_31__bench === 1'bx)) begin
				n3_odata_p0_31__flag <= 1'b1;
			end else begin
				n3_odata_p0_31__flag<= 1'b0;
			end
			if(!(n3_odata_p0_32__gfpga === n3_odata_p0_32__bench) && !(n3_odata_p0_32__bench === 1'bx)) begin
				n3_odata_p0_32__flag <= 1'b1;
			end else begin
				n3_odata_p0_32__flag<= 1'b0;
			end
			if(!(n3_odata_p0_33__gfpga === n3_odata_p0_33__bench) && !(n3_odata_p0_33__bench === 1'bx)) begin
				n3_odata_p0_33__flag <= 1'b1;
			end else begin
				n3_odata_p0_33__flag<= 1'b0;
			end
			if(!(n3_odata_p0_34__gfpga === n3_odata_p0_34__bench) && !(n3_odata_p0_34__bench === 1'bx)) begin
				n3_odata_p0_34__flag <= 1'b1;
			end else begin
				n3_odata_p0_34__flag<= 1'b0;
			end
			if(!(n3_ovalid_p0_gfpga === n3_ovalid_p0_bench) && !(n3_ovalid_p0_bench === 1'bx)) begin
				n3_ovalid_p0_flag <= 1'b1;
			end else begin
				n3_ovalid_p0_flag<= 1'b0;
			end
			if(!(n4_ordy_p0_0__gfpga === n4_ordy_p0_0__bench) && !(n4_ordy_p0_0__bench === 1'bx)) begin
				n4_ordy_p0_0__flag <= 1'b1;
			end else begin
				n4_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n4_ordy_p0_1__gfpga === n4_ordy_p0_1__bench) && !(n4_ordy_p0_1__bench === 1'bx)) begin
				n4_ordy_p0_1__flag <= 1'b1;
			end else begin
				n4_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n4_odata_p0_0__gfpga === n4_odata_p0_0__bench) && !(n4_odata_p0_0__bench === 1'bx)) begin
				n4_odata_p0_0__flag <= 1'b1;
			end else begin
				n4_odata_p0_0__flag<= 1'b0;
			end
			if(!(n4_odata_p0_1__gfpga === n4_odata_p0_1__bench) && !(n4_odata_p0_1__bench === 1'bx)) begin
				n4_odata_p0_1__flag <= 1'b1;
			end else begin
				n4_odata_p0_1__flag<= 1'b0;
			end
			if(!(n4_odata_p0_2__gfpga === n4_odata_p0_2__bench) && !(n4_odata_p0_2__bench === 1'bx)) begin
				n4_odata_p0_2__flag <= 1'b1;
			end else begin
				n4_odata_p0_2__flag<= 1'b0;
			end
			if(!(n4_odata_p0_3__gfpga === n4_odata_p0_3__bench) && !(n4_odata_p0_3__bench === 1'bx)) begin
				n4_odata_p0_3__flag <= 1'b1;
			end else begin
				n4_odata_p0_3__flag<= 1'b0;
			end
			if(!(n4_odata_p0_4__gfpga === n4_odata_p0_4__bench) && !(n4_odata_p0_4__bench === 1'bx)) begin
				n4_odata_p0_4__flag <= 1'b1;
			end else begin
				n4_odata_p0_4__flag<= 1'b0;
			end
			if(!(n4_odata_p0_5__gfpga === n4_odata_p0_5__bench) && !(n4_odata_p0_5__bench === 1'bx)) begin
				n4_odata_p0_5__flag <= 1'b1;
			end else begin
				n4_odata_p0_5__flag<= 1'b0;
			end
			if(!(n4_odata_p0_6__gfpga === n4_odata_p0_6__bench) && !(n4_odata_p0_6__bench === 1'bx)) begin
				n4_odata_p0_6__flag <= 1'b1;
			end else begin
				n4_odata_p0_6__flag<= 1'b0;
			end
			if(!(n4_odata_p0_7__gfpga === n4_odata_p0_7__bench) && !(n4_odata_p0_7__bench === 1'bx)) begin
				n4_odata_p0_7__flag <= 1'b1;
			end else begin
				n4_odata_p0_7__flag<= 1'b0;
			end
			if(!(n4_odata_p0_8__gfpga === n4_odata_p0_8__bench) && !(n4_odata_p0_8__bench === 1'bx)) begin
				n4_odata_p0_8__flag <= 1'b1;
			end else begin
				n4_odata_p0_8__flag<= 1'b0;
			end
			if(!(n4_odata_p0_9__gfpga === n4_odata_p0_9__bench) && !(n4_odata_p0_9__bench === 1'bx)) begin
				n4_odata_p0_9__flag <= 1'b1;
			end else begin
				n4_odata_p0_9__flag<= 1'b0;
			end
			if(!(n4_odata_p0_10__gfpga === n4_odata_p0_10__bench) && !(n4_odata_p0_10__bench === 1'bx)) begin
				n4_odata_p0_10__flag <= 1'b1;
			end else begin
				n4_odata_p0_10__flag<= 1'b0;
			end
			if(!(n4_odata_p0_11__gfpga === n4_odata_p0_11__bench) && !(n4_odata_p0_11__bench === 1'bx)) begin
				n4_odata_p0_11__flag <= 1'b1;
			end else begin
				n4_odata_p0_11__flag<= 1'b0;
			end
			if(!(n4_odata_p0_12__gfpga === n4_odata_p0_12__bench) && !(n4_odata_p0_12__bench === 1'bx)) begin
				n4_odata_p0_12__flag <= 1'b1;
			end else begin
				n4_odata_p0_12__flag<= 1'b0;
			end
			if(!(n4_odata_p0_13__gfpga === n4_odata_p0_13__bench) && !(n4_odata_p0_13__bench === 1'bx)) begin
				n4_odata_p0_13__flag <= 1'b1;
			end else begin
				n4_odata_p0_13__flag<= 1'b0;
			end
			if(!(n4_odata_p0_14__gfpga === n4_odata_p0_14__bench) && !(n4_odata_p0_14__bench === 1'bx)) begin
				n4_odata_p0_14__flag <= 1'b1;
			end else begin
				n4_odata_p0_14__flag<= 1'b0;
			end
			if(!(n4_odata_p0_15__gfpga === n4_odata_p0_15__bench) && !(n4_odata_p0_15__bench === 1'bx)) begin
				n4_odata_p0_15__flag <= 1'b1;
			end else begin
				n4_odata_p0_15__flag<= 1'b0;
			end
			if(!(n4_odata_p0_16__gfpga === n4_odata_p0_16__bench) && !(n4_odata_p0_16__bench === 1'bx)) begin
				n4_odata_p0_16__flag <= 1'b1;
			end else begin
				n4_odata_p0_16__flag<= 1'b0;
			end
			if(!(n4_odata_p0_17__gfpga === n4_odata_p0_17__bench) && !(n4_odata_p0_17__bench === 1'bx)) begin
				n4_odata_p0_17__flag <= 1'b1;
			end else begin
				n4_odata_p0_17__flag<= 1'b0;
			end
			if(!(n4_odata_p0_18__gfpga === n4_odata_p0_18__bench) && !(n4_odata_p0_18__bench === 1'bx)) begin
				n4_odata_p0_18__flag <= 1'b1;
			end else begin
				n4_odata_p0_18__flag<= 1'b0;
			end
			if(!(n4_odata_p0_19__gfpga === n4_odata_p0_19__bench) && !(n4_odata_p0_19__bench === 1'bx)) begin
				n4_odata_p0_19__flag <= 1'b1;
			end else begin
				n4_odata_p0_19__flag<= 1'b0;
			end
			if(!(n4_odata_p0_20__gfpga === n4_odata_p0_20__bench) && !(n4_odata_p0_20__bench === 1'bx)) begin
				n4_odata_p0_20__flag <= 1'b1;
			end else begin
				n4_odata_p0_20__flag<= 1'b0;
			end
			if(!(n4_odata_p0_21__gfpga === n4_odata_p0_21__bench) && !(n4_odata_p0_21__bench === 1'bx)) begin
				n4_odata_p0_21__flag <= 1'b1;
			end else begin
				n4_odata_p0_21__flag<= 1'b0;
			end
			if(!(n4_odata_p0_22__gfpga === n4_odata_p0_22__bench) && !(n4_odata_p0_22__bench === 1'bx)) begin
				n4_odata_p0_22__flag <= 1'b1;
			end else begin
				n4_odata_p0_22__flag<= 1'b0;
			end
			if(!(n4_odata_p0_23__gfpga === n4_odata_p0_23__bench) && !(n4_odata_p0_23__bench === 1'bx)) begin
				n4_odata_p0_23__flag <= 1'b1;
			end else begin
				n4_odata_p0_23__flag<= 1'b0;
			end
			if(!(n4_odata_p0_24__gfpga === n4_odata_p0_24__bench) && !(n4_odata_p0_24__bench === 1'bx)) begin
				n4_odata_p0_24__flag <= 1'b1;
			end else begin
				n4_odata_p0_24__flag<= 1'b0;
			end
			if(!(n4_odata_p0_25__gfpga === n4_odata_p0_25__bench) && !(n4_odata_p0_25__bench === 1'bx)) begin
				n4_odata_p0_25__flag <= 1'b1;
			end else begin
				n4_odata_p0_25__flag<= 1'b0;
			end
			if(!(n4_odata_p0_26__gfpga === n4_odata_p0_26__bench) && !(n4_odata_p0_26__bench === 1'bx)) begin
				n4_odata_p0_26__flag <= 1'b1;
			end else begin
				n4_odata_p0_26__flag<= 1'b0;
			end
			if(!(n4_odata_p0_27__gfpga === n4_odata_p0_27__bench) && !(n4_odata_p0_27__bench === 1'bx)) begin
				n4_odata_p0_27__flag <= 1'b1;
			end else begin
				n4_odata_p0_27__flag<= 1'b0;
			end
			if(!(n4_odata_p0_28__gfpga === n4_odata_p0_28__bench) && !(n4_odata_p0_28__bench === 1'bx)) begin
				n4_odata_p0_28__flag <= 1'b1;
			end else begin
				n4_odata_p0_28__flag<= 1'b0;
			end
			if(!(n4_odata_p0_29__gfpga === n4_odata_p0_29__bench) && !(n4_odata_p0_29__bench === 1'bx)) begin
				n4_odata_p0_29__flag <= 1'b1;
			end else begin
				n4_odata_p0_29__flag<= 1'b0;
			end
			if(!(n4_odata_p0_30__gfpga === n4_odata_p0_30__bench) && !(n4_odata_p0_30__bench === 1'bx)) begin
				n4_odata_p0_30__flag <= 1'b1;
			end else begin
				n4_odata_p0_30__flag<= 1'b0;
			end
			if(!(n4_odata_p0_31__gfpga === n4_odata_p0_31__bench) && !(n4_odata_p0_31__bench === 1'bx)) begin
				n4_odata_p0_31__flag <= 1'b1;
			end else begin
				n4_odata_p0_31__flag<= 1'b0;
			end
			if(!(n4_odata_p0_32__gfpga === n4_odata_p0_32__bench) && !(n4_odata_p0_32__bench === 1'bx)) begin
				n4_odata_p0_32__flag <= 1'b1;
			end else begin
				n4_odata_p0_32__flag<= 1'b0;
			end
			if(!(n4_odata_p0_33__gfpga === n4_odata_p0_33__bench) && !(n4_odata_p0_33__bench === 1'bx)) begin
				n4_odata_p0_33__flag <= 1'b1;
			end else begin
				n4_odata_p0_33__flag<= 1'b0;
			end
			if(!(n4_odata_p0_34__gfpga === n4_odata_p0_34__bench) && !(n4_odata_p0_34__bench === 1'bx)) begin
				n4_odata_p0_34__flag <= 1'b1;
			end else begin
				n4_odata_p0_34__flag<= 1'b0;
			end
			if(!(n4_ovalid_p0_gfpga === n4_ovalid_p0_bench) && !(n4_ovalid_p0_bench === 1'bx)) begin
				n4_ovalid_p0_flag <= 1'b1;
			end else begin
				n4_ovalid_p0_flag<= 1'b0;
			end
			if(!(n5_ordy_p0_0__gfpga === n5_ordy_p0_0__bench) && !(n5_ordy_p0_0__bench === 1'bx)) begin
				n5_ordy_p0_0__flag <= 1'b1;
			end else begin
				n5_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n5_ordy_p0_1__gfpga === n5_ordy_p0_1__bench) && !(n5_ordy_p0_1__bench === 1'bx)) begin
				n5_ordy_p0_1__flag <= 1'b1;
			end else begin
				n5_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n5_odata_p0_0__gfpga === n5_odata_p0_0__bench) && !(n5_odata_p0_0__bench === 1'bx)) begin
				n5_odata_p0_0__flag <= 1'b1;
			end else begin
				n5_odata_p0_0__flag<= 1'b0;
			end
			if(!(n5_odata_p0_1__gfpga === n5_odata_p0_1__bench) && !(n5_odata_p0_1__bench === 1'bx)) begin
				n5_odata_p0_1__flag <= 1'b1;
			end else begin
				n5_odata_p0_1__flag<= 1'b0;
			end
			if(!(n5_odata_p0_2__gfpga === n5_odata_p0_2__bench) && !(n5_odata_p0_2__bench === 1'bx)) begin
				n5_odata_p0_2__flag <= 1'b1;
			end else begin
				n5_odata_p0_2__flag<= 1'b0;
			end
			if(!(n5_odata_p0_3__gfpga === n5_odata_p0_3__bench) && !(n5_odata_p0_3__bench === 1'bx)) begin
				n5_odata_p0_3__flag <= 1'b1;
			end else begin
				n5_odata_p0_3__flag<= 1'b0;
			end
			if(!(n5_odata_p0_4__gfpga === n5_odata_p0_4__bench) && !(n5_odata_p0_4__bench === 1'bx)) begin
				n5_odata_p0_4__flag <= 1'b1;
			end else begin
				n5_odata_p0_4__flag<= 1'b0;
			end
			if(!(n5_odata_p0_5__gfpga === n5_odata_p0_5__bench) && !(n5_odata_p0_5__bench === 1'bx)) begin
				n5_odata_p0_5__flag <= 1'b1;
			end else begin
				n5_odata_p0_5__flag<= 1'b0;
			end
			if(!(n5_odata_p0_6__gfpga === n5_odata_p0_6__bench) && !(n5_odata_p0_6__bench === 1'bx)) begin
				n5_odata_p0_6__flag <= 1'b1;
			end else begin
				n5_odata_p0_6__flag<= 1'b0;
			end
			if(!(n5_odata_p0_7__gfpga === n5_odata_p0_7__bench) && !(n5_odata_p0_7__bench === 1'bx)) begin
				n5_odata_p0_7__flag <= 1'b1;
			end else begin
				n5_odata_p0_7__flag<= 1'b0;
			end
			if(!(n5_odata_p0_8__gfpga === n5_odata_p0_8__bench) && !(n5_odata_p0_8__bench === 1'bx)) begin
				n5_odata_p0_8__flag <= 1'b1;
			end else begin
				n5_odata_p0_8__flag<= 1'b0;
			end
			if(!(n5_odata_p0_9__gfpga === n5_odata_p0_9__bench) && !(n5_odata_p0_9__bench === 1'bx)) begin
				n5_odata_p0_9__flag <= 1'b1;
			end else begin
				n5_odata_p0_9__flag<= 1'b0;
			end
			if(!(n5_odata_p0_10__gfpga === n5_odata_p0_10__bench) && !(n5_odata_p0_10__bench === 1'bx)) begin
				n5_odata_p0_10__flag <= 1'b1;
			end else begin
				n5_odata_p0_10__flag<= 1'b0;
			end
			if(!(n5_odata_p0_11__gfpga === n5_odata_p0_11__bench) && !(n5_odata_p0_11__bench === 1'bx)) begin
				n5_odata_p0_11__flag <= 1'b1;
			end else begin
				n5_odata_p0_11__flag<= 1'b0;
			end
			if(!(n5_odata_p0_12__gfpga === n5_odata_p0_12__bench) && !(n5_odata_p0_12__bench === 1'bx)) begin
				n5_odata_p0_12__flag <= 1'b1;
			end else begin
				n5_odata_p0_12__flag<= 1'b0;
			end
			if(!(n5_odata_p0_13__gfpga === n5_odata_p0_13__bench) && !(n5_odata_p0_13__bench === 1'bx)) begin
				n5_odata_p0_13__flag <= 1'b1;
			end else begin
				n5_odata_p0_13__flag<= 1'b0;
			end
			if(!(n5_odata_p0_14__gfpga === n5_odata_p0_14__bench) && !(n5_odata_p0_14__bench === 1'bx)) begin
				n5_odata_p0_14__flag <= 1'b1;
			end else begin
				n5_odata_p0_14__flag<= 1'b0;
			end
			if(!(n5_odata_p0_15__gfpga === n5_odata_p0_15__bench) && !(n5_odata_p0_15__bench === 1'bx)) begin
				n5_odata_p0_15__flag <= 1'b1;
			end else begin
				n5_odata_p0_15__flag<= 1'b0;
			end
			if(!(n5_odata_p0_16__gfpga === n5_odata_p0_16__bench) && !(n5_odata_p0_16__bench === 1'bx)) begin
				n5_odata_p0_16__flag <= 1'b1;
			end else begin
				n5_odata_p0_16__flag<= 1'b0;
			end
			if(!(n5_odata_p0_17__gfpga === n5_odata_p0_17__bench) && !(n5_odata_p0_17__bench === 1'bx)) begin
				n5_odata_p0_17__flag <= 1'b1;
			end else begin
				n5_odata_p0_17__flag<= 1'b0;
			end
			if(!(n5_odata_p0_18__gfpga === n5_odata_p0_18__bench) && !(n5_odata_p0_18__bench === 1'bx)) begin
				n5_odata_p0_18__flag <= 1'b1;
			end else begin
				n5_odata_p0_18__flag<= 1'b0;
			end
			if(!(n5_odata_p0_19__gfpga === n5_odata_p0_19__bench) && !(n5_odata_p0_19__bench === 1'bx)) begin
				n5_odata_p0_19__flag <= 1'b1;
			end else begin
				n5_odata_p0_19__flag<= 1'b0;
			end
			if(!(n5_odata_p0_20__gfpga === n5_odata_p0_20__bench) && !(n5_odata_p0_20__bench === 1'bx)) begin
				n5_odata_p0_20__flag <= 1'b1;
			end else begin
				n5_odata_p0_20__flag<= 1'b0;
			end
			if(!(n5_odata_p0_21__gfpga === n5_odata_p0_21__bench) && !(n5_odata_p0_21__bench === 1'bx)) begin
				n5_odata_p0_21__flag <= 1'b1;
			end else begin
				n5_odata_p0_21__flag<= 1'b0;
			end
			if(!(n5_odata_p0_22__gfpga === n5_odata_p0_22__bench) && !(n5_odata_p0_22__bench === 1'bx)) begin
				n5_odata_p0_22__flag <= 1'b1;
			end else begin
				n5_odata_p0_22__flag<= 1'b0;
			end
			if(!(n5_odata_p0_23__gfpga === n5_odata_p0_23__bench) && !(n5_odata_p0_23__bench === 1'bx)) begin
				n5_odata_p0_23__flag <= 1'b1;
			end else begin
				n5_odata_p0_23__flag<= 1'b0;
			end
			if(!(n5_odata_p0_24__gfpga === n5_odata_p0_24__bench) && !(n5_odata_p0_24__bench === 1'bx)) begin
				n5_odata_p0_24__flag <= 1'b1;
			end else begin
				n5_odata_p0_24__flag<= 1'b0;
			end
			if(!(n5_odata_p0_25__gfpga === n5_odata_p0_25__bench) && !(n5_odata_p0_25__bench === 1'bx)) begin
				n5_odata_p0_25__flag <= 1'b1;
			end else begin
				n5_odata_p0_25__flag<= 1'b0;
			end
			if(!(n5_odata_p0_26__gfpga === n5_odata_p0_26__bench) && !(n5_odata_p0_26__bench === 1'bx)) begin
				n5_odata_p0_26__flag <= 1'b1;
			end else begin
				n5_odata_p0_26__flag<= 1'b0;
			end
			if(!(n5_odata_p0_27__gfpga === n5_odata_p0_27__bench) && !(n5_odata_p0_27__bench === 1'bx)) begin
				n5_odata_p0_27__flag <= 1'b1;
			end else begin
				n5_odata_p0_27__flag<= 1'b0;
			end
			if(!(n5_odata_p0_28__gfpga === n5_odata_p0_28__bench) && !(n5_odata_p0_28__bench === 1'bx)) begin
				n5_odata_p0_28__flag <= 1'b1;
			end else begin
				n5_odata_p0_28__flag<= 1'b0;
			end
			if(!(n5_odata_p0_29__gfpga === n5_odata_p0_29__bench) && !(n5_odata_p0_29__bench === 1'bx)) begin
				n5_odata_p0_29__flag <= 1'b1;
			end else begin
				n5_odata_p0_29__flag<= 1'b0;
			end
			if(!(n5_odata_p0_30__gfpga === n5_odata_p0_30__bench) && !(n5_odata_p0_30__bench === 1'bx)) begin
				n5_odata_p0_30__flag <= 1'b1;
			end else begin
				n5_odata_p0_30__flag<= 1'b0;
			end
			if(!(n5_odata_p0_31__gfpga === n5_odata_p0_31__bench) && !(n5_odata_p0_31__bench === 1'bx)) begin
				n5_odata_p0_31__flag <= 1'b1;
			end else begin
				n5_odata_p0_31__flag<= 1'b0;
			end
			if(!(n5_odata_p0_32__gfpga === n5_odata_p0_32__bench) && !(n5_odata_p0_32__bench === 1'bx)) begin
				n5_odata_p0_32__flag <= 1'b1;
			end else begin
				n5_odata_p0_32__flag<= 1'b0;
			end
			if(!(n5_odata_p0_33__gfpga === n5_odata_p0_33__bench) && !(n5_odata_p0_33__bench === 1'bx)) begin
				n5_odata_p0_33__flag <= 1'b1;
			end else begin
				n5_odata_p0_33__flag<= 1'b0;
			end
			if(!(n5_odata_p0_34__gfpga === n5_odata_p0_34__bench) && !(n5_odata_p0_34__bench === 1'bx)) begin
				n5_odata_p0_34__flag <= 1'b1;
			end else begin
				n5_odata_p0_34__flag<= 1'b0;
			end
			if(!(n5_ovalid_p0_gfpga === n5_ovalid_p0_bench) && !(n5_ovalid_p0_bench === 1'bx)) begin
				n5_ovalid_p0_flag <= 1'b1;
			end else begin
				n5_ovalid_p0_flag<= 1'b0;
			end
			if(!(n6_ordy_p0_0__gfpga === n6_ordy_p0_0__bench) && !(n6_ordy_p0_0__bench === 1'bx)) begin
				n6_ordy_p0_0__flag <= 1'b1;
			end else begin
				n6_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n6_ordy_p0_1__gfpga === n6_ordy_p0_1__bench) && !(n6_ordy_p0_1__bench === 1'bx)) begin
				n6_ordy_p0_1__flag <= 1'b1;
			end else begin
				n6_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n6_odata_p0_0__gfpga === n6_odata_p0_0__bench) && !(n6_odata_p0_0__bench === 1'bx)) begin
				n6_odata_p0_0__flag <= 1'b1;
			end else begin
				n6_odata_p0_0__flag<= 1'b0;
			end
			if(!(n6_odata_p0_1__gfpga === n6_odata_p0_1__bench) && !(n6_odata_p0_1__bench === 1'bx)) begin
				n6_odata_p0_1__flag <= 1'b1;
			end else begin
				n6_odata_p0_1__flag<= 1'b0;
			end
			if(!(n6_odata_p0_2__gfpga === n6_odata_p0_2__bench) && !(n6_odata_p0_2__bench === 1'bx)) begin
				n6_odata_p0_2__flag <= 1'b1;
			end else begin
				n6_odata_p0_2__flag<= 1'b0;
			end
			if(!(n6_odata_p0_3__gfpga === n6_odata_p0_3__bench) && !(n6_odata_p0_3__bench === 1'bx)) begin
				n6_odata_p0_3__flag <= 1'b1;
			end else begin
				n6_odata_p0_3__flag<= 1'b0;
			end
			if(!(n6_odata_p0_4__gfpga === n6_odata_p0_4__bench) && !(n6_odata_p0_4__bench === 1'bx)) begin
				n6_odata_p0_4__flag <= 1'b1;
			end else begin
				n6_odata_p0_4__flag<= 1'b0;
			end
			if(!(n6_odata_p0_5__gfpga === n6_odata_p0_5__bench) && !(n6_odata_p0_5__bench === 1'bx)) begin
				n6_odata_p0_5__flag <= 1'b1;
			end else begin
				n6_odata_p0_5__flag<= 1'b0;
			end
			if(!(n6_odata_p0_6__gfpga === n6_odata_p0_6__bench) && !(n6_odata_p0_6__bench === 1'bx)) begin
				n6_odata_p0_6__flag <= 1'b1;
			end else begin
				n6_odata_p0_6__flag<= 1'b0;
			end
			if(!(n6_odata_p0_7__gfpga === n6_odata_p0_7__bench) && !(n6_odata_p0_7__bench === 1'bx)) begin
				n6_odata_p0_7__flag <= 1'b1;
			end else begin
				n6_odata_p0_7__flag<= 1'b0;
			end
			if(!(n6_odata_p0_8__gfpga === n6_odata_p0_8__bench) && !(n6_odata_p0_8__bench === 1'bx)) begin
				n6_odata_p0_8__flag <= 1'b1;
			end else begin
				n6_odata_p0_8__flag<= 1'b0;
			end
			if(!(n6_odata_p0_9__gfpga === n6_odata_p0_9__bench) && !(n6_odata_p0_9__bench === 1'bx)) begin
				n6_odata_p0_9__flag <= 1'b1;
			end else begin
				n6_odata_p0_9__flag<= 1'b0;
			end
			if(!(n6_odata_p0_10__gfpga === n6_odata_p0_10__bench) && !(n6_odata_p0_10__bench === 1'bx)) begin
				n6_odata_p0_10__flag <= 1'b1;
			end else begin
				n6_odata_p0_10__flag<= 1'b0;
			end
			if(!(n6_odata_p0_11__gfpga === n6_odata_p0_11__bench) && !(n6_odata_p0_11__bench === 1'bx)) begin
				n6_odata_p0_11__flag <= 1'b1;
			end else begin
				n6_odata_p0_11__flag<= 1'b0;
			end
			if(!(n6_odata_p0_12__gfpga === n6_odata_p0_12__bench) && !(n6_odata_p0_12__bench === 1'bx)) begin
				n6_odata_p0_12__flag <= 1'b1;
			end else begin
				n6_odata_p0_12__flag<= 1'b0;
			end
			if(!(n6_odata_p0_13__gfpga === n6_odata_p0_13__bench) && !(n6_odata_p0_13__bench === 1'bx)) begin
				n6_odata_p0_13__flag <= 1'b1;
			end else begin
				n6_odata_p0_13__flag<= 1'b0;
			end
			if(!(n6_odata_p0_14__gfpga === n6_odata_p0_14__bench) && !(n6_odata_p0_14__bench === 1'bx)) begin
				n6_odata_p0_14__flag <= 1'b1;
			end else begin
				n6_odata_p0_14__flag<= 1'b0;
			end
			if(!(n6_odata_p0_15__gfpga === n6_odata_p0_15__bench) && !(n6_odata_p0_15__bench === 1'bx)) begin
				n6_odata_p0_15__flag <= 1'b1;
			end else begin
				n6_odata_p0_15__flag<= 1'b0;
			end
			if(!(n6_odata_p0_16__gfpga === n6_odata_p0_16__bench) && !(n6_odata_p0_16__bench === 1'bx)) begin
				n6_odata_p0_16__flag <= 1'b1;
			end else begin
				n6_odata_p0_16__flag<= 1'b0;
			end
			if(!(n6_odata_p0_17__gfpga === n6_odata_p0_17__bench) && !(n6_odata_p0_17__bench === 1'bx)) begin
				n6_odata_p0_17__flag <= 1'b1;
			end else begin
				n6_odata_p0_17__flag<= 1'b0;
			end
			if(!(n6_odata_p0_18__gfpga === n6_odata_p0_18__bench) && !(n6_odata_p0_18__bench === 1'bx)) begin
				n6_odata_p0_18__flag <= 1'b1;
			end else begin
				n6_odata_p0_18__flag<= 1'b0;
			end
			if(!(n6_odata_p0_19__gfpga === n6_odata_p0_19__bench) && !(n6_odata_p0_19__bench === 1'bx)) begin
				n6_odata_p0_19__flag <= 1'b1;
			end else begin
				n6_odata_p0_19__flag<= 1'b0;
			end
			if(!(n6_odata_p0_20__gfpga === n6_odata_p0_20__bench) && !(n6_odata_p0_20__bench === 1'bx)) begin
				n6_odata_p0_20__flag <= 1'b1;
			end else begin
				n6_odata_p0_20__flag<= 1'b0;
			end
			if(!(n6_odata_p0_21__gfpga === n6_odata_p0_21__bench) && !(n6_odata_p0_21__bench === 1'bx)) begin
				n6_odata_p0_21__flag <= 1'b1;
			end else begin
				n6_odata_p0_21__flag<= 1'b0;
			end
			if(!(n6_odata_p0_22__gfpga === n6_odata_p0_22__bench) && !(n6_odata_p0_22__bench === 1'bx)) begin
				n6_odata_p0_22__flag <= 1'b1;
			end else begin
				n6_odata_p0_22__flag<= 1'b0;
			end
			if(!(n6_odata_p0_23__gfpga === n6_odata_p0_23__bench) && !(n6_odata_p0_23__bench === 1'bx)) begin
				n6_odata_p0_23__flag <= 1'b1;
			end else begin
				n6_odata_p0_23__flag<= 1'b0;
			end
			if(!(n6_odata_p0_24__gfpga === n6_odata_p0_24__bench) && !(n6_odata_p0_24__bench === 1'bx)) begin
				n6_odata_p0_24__flag <= 1'b1;
			end else begin
				n6_odata_p0_24__flag<= 1'b0;
			end
			if(!(n6_odata_p0_25__gfpga === n6_odata_p0_25__bench) && !(n6_odata_p0_25__bench === 1'bx)) begin
				n6_odata_p0_25__flag <= 1'b1;
			end else begin
				n6_odata_p0_25__flag<= 1'b0;
			end
			if(!(n6_odata_p0_26__gfpga === n6_odata_p0_26__bench) && !(n6_odata_p0_26__bench === 1'bx)) begin
				n6_odata_p0_26__flag <= 1'b1;
			end else begin
				n6_odata_p0_26__flag<= 1'b0;
			end
			if(!(n6_odata_p0_27__gfpga === n6_odata_p0_27__bench) && !(n6_odata_p0_27__bench === 1'bx)) begin
				n6_odata_p0_27__flag <= 1'b1;
			end else begin
				n6_odata_p0_27__flag<= 1'b0;
			end
			if(!(n6_odata_p0_28__gfpga === n6_odata_p0_28__bench) && !(n6_odata_p0_28__bench === 1'bx)) begin
				n6_odata_p0_28__flag <= 1'b1;
			end else begin
				n6_odata_p0_28__flag<= 1'b0;
			end
			if(!(n6_odata_p0_29__gfpga === n6_odata_p0_29__bench) && !(n6_odata_p0_29__bench === 1'bx)) begin
				n6_odata_p0_29__flag <= 1'b1;
			end else begin
				n6_odata_p0_29__flag<= 1'b0;
			end
			if(!(n6_odata_p0_30__gfpga === n6_odata_p0_30__bench) && !(n6_odata_p0_30__bench === 1'bx)) begin
				n6_odata_p0_30__flag <= 1'b1;
			end else begin
				n6_odata_p0_30__flag<= 1'b0;
			end
			if(!(n6_odata_p0_31__gfpga === n6_odata_p0_31__bench) && !(n6_odata_p0_31__bench === 1'bx)) begin
				n6_odata_p0_31__flag <= 1'b1;
			end else begin
				n6_odata_p0_31__flag<= 1'b0;
			end
			if(!(n6_odata_p0_32__gfpga === n6_odata_p0_32__bench) && !(n6_odata_p0_32__bench === 1'bx)) begin
				n6_odata_p0_32__flag <= 1'b1;
			end else begin
				n6_odata_p0_32__flag<= 1'b0;
			end
			if(!(n6_odata_p0_33__gfpga === n6_odata_p0_33__bench) && !(n6_odata_p0_33__bench === 1'bx)) begin
				n6_odata_p0_33__flag <= 1'b1;
			end else begin
				n6_odata_p0_33__flag<= 1'b0;
			end
			if(!(n6_odata_p0_34__gfpga === n6_odata_p0_34__bench) && !(n6_odata_p0_34__bench === 1'bx)) begin
				n6_odata_p0_34__flag <= 1'b1;
			end else begin
				n6_odata_p0_34__flag<= 1'b0;
			end
			if(!(n6_ovalid_p0_gfpga === n6_ovalid_p0_bench) && !(n6_ovalid_p0_bench === 1'bx)) begin
				n6_ovalid_p0_flag <= 1'b1;
			end else begin
				n6_ovalid_p0_flag<= 1'b0;
			end
			if(!(n7_ordy_p0_0__gfpga === n7_ordy_p0_0__bench) && !(n7_ordy_p0_0__bench === 1'bx)) begin
				n7_ordy_p0_0__flag <= 1'b1;
			end else begin
				n7_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n7_ordy_p0_1__gfpga === n7_ordy_p0_1__bench) && !(n7_ordy_p0_1__bench === 1'bx)) begin
				n7_ordy_p0_1__flag <= 1'b1;
			end else begin
				n7_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n7_odata_p0_0__gfpga === n7_odata_p0_0__bench) && !(n7_odata_p0_0__bench === 1'bx)) begin
				n7_odata_p0_0__flag <= 1'b1;
			end else begin
				n7_odata_p0_0__flag<= 1'b0;
			end
			if(!(n7_odata_p0_1__gfpga === n7_odata_p0_1__bench) && !(n7_odata_p0_1__bench === 1'bx)) begin
				n7_odata_p0_1__flag <= 1'b1;
			end else begin
				n7_odata_p0_1__flag<= 1'b0;
			end
			if(!(n7_odata_p0_2__gfpga === n7_odata_p0_2__bench) && !(n7_odata_p0_2__bench === 1'bx)) begin
				n7_odata_p0_2__flag <= 1'b1;
			end else begin
				n7_odata_p0_2__flag<= 1'b0;
			end
			if(!(n7_odata_p0_3__gfpga === n7_odata_p0_3__bench) && !(n7_odata_p0_3__bench === 1'bx)) begin
				n7_odata_p0_3__flag <= 1'b1;
			end else begin
				n7_odata_p0_3__flag<= 1'b0;
			end
			if(!(n7_odata_p0_4__gfpga === n7_odata_p0_4__bench) && !(n7_odata_p0_4__bench === 1'bx)) begin
				n7_odata_p0_4__flag <= 1'b1;
			end else begin
				n7_odata_p0_4__flag<= 1'b0;
			end
			if(!(n7_odata_p0_5__gfpga === n7_odata_p0_5__bench) && !(n7_odata_p0_5__bench === 1'bx)) begin
				n7_odata_p0_5__flag <= 1'b1;
			end else begin
				n7_odata_p0_5__flag<= 1'b0;
			end
			if(!(n7_odata_p0_6__gfpga === n7_odata_p0_6__bench) && !(n7_odata_p0_6__bench === 1'bx)) begin
				n7_odata_p0_6__flag <= 1'b1;
			end else begin
				n7_odata_p0_6__flag<= 1'b0;
			end
			if(!(n7_odata_p0_7__gfpga === n7_odata_p0_7__bench) && !(n7_odata_p0_7__bench === 1'bx)) begin
				n7_odata_p0_7__flag <= 1'b1;
			end else begin
				n7_odata_p0_7__flag<= 1'b0;
			end
			if(!(n7_odata_p0_8__gfpga === n7_odata_p0_8__bench) && !(n7_odata_p0_8__bench === 1'bx)) begin
				n7_odata_p0_8__flag <= 1'b1;
			end else begin
				n7_odata_p0_8__flag<= 1'b0;
			end
			if(!(n7_odata_p0_9__gfpga === n7_odata_p0_9__bench) && !(n7_odata_p0_9__bench === 1'bx)) begin
				n7_odata_p0_9__flag <= 1'b1;
			end else begin
				n7_odata_p0_9__flag<= 1'b0;
			end
			if(!(n7_odata_p0_10__gfpga === n7_odata_p0_10__bench) && !(n7_odata_p0_10__bench === 1'bx)) begin
				n7_odata_p0_10__flag <= 1'b1;
			end else begin
				n7_odata_p0_10__flag<= 1'b0;
			end
			if(!(n7_odata_p0_11__gfpga === n7_odata_p0_11__bench) && !(n7_odata_p0_11__bench === 1'bx)) begin
				n7_odata_p0_11__flag <= 1'b1;
			end else begin
				n7_odata_p0_11__flag<= 1'b0;
			end
			if(!(n7_odata_p0_12__gfpga === n7_odata_p0_12__bench) && !(n7_odata_p0_12__bench === 1'bx)) begin
				n7_odata_p0_12__flag <= 1'b1;
			end else begin
				n7_odata_p0_12__flag<= 1'b0;
			end
			if(!(n7_odata_p0_13__gfpga === n7_odata_p0_13__bench) && !(n7_odata_p0_13__bench === 1'bx)) begin
				n7_odata_p0_13__flag <= 1'b1;
			end else begin
				n7_odata_p0_13__flag<= 1'b0;
			end
			if(!(n7_odata_p0_14__gfpga === n7_odata_p0_14__bench) && !(n7_odata_p0_14__bench === 1'bx)) begin
				n7_odata_p0_14__flag <= 1'b1;
			end else begin
				n7_odata_p0_14__flag<= 1'b0;
			end
			if(!(n7_odata_p0_15__gfpga === n7_odata_p0_15__bench) && !(n7_odata_p0_15__bench === 1'bx)) begin
				n7_odata_p0_15__flag <= 1'b1;
			end else begin
				n7_odata_p0_15__flag<= 1'b0;
			end
			if(!(n7_odata_p0_16__gfpga === n7_odata_p0_16__bench) && !(n7_odata_p0_16__bench === 1'bx)) begin
				n7_odata_p0_16__flag <= 1'b1;
			end else begin
				n7_odata_p0_16__flag<= 1'b0;
			end
			if(!(n7_odata_p0_17__gfpga === n7_odata_p0_17__bench) && !(n7_odata_p0_17__bench === 1'bx)) begin
				n7_odata_p0_17__flag <= 1'b1;
			end else begin
				n7_odata_p0_17__flag<= 1'b0;
			end
			if(!(n7_odata_p0_18__gfpga === n7_odata_p0_18__bench) && !(n7_odata_p0_18__bench === 1'bx)) begin
				n7_odata_p0_18__flag <= 1'b1;
			end else begin
				n7_odata_p0_18__flag<= 1'b0;
			end
			if(!(n7_odata_p0_19__gfpga === n7_odata_p0_19__bench) && !(n7_odata_p0_19__bench === 1'bx)) begin
				n7_odata_p0_19__flag <= 1'b1;
			end else begin
				n7_odata_p0_19__flag<= 1'b0;
			end
			if(!(n7_odata_p0_20__gfpga === n7_odata_p0_20__bench) && !(n7_odata_p0_20__bench === 1'bx)) begin
				n7_odata_p0_20__flag <= 1'b1;
			end else begin
				n7_odata_p0_20__flag<= 1'b0;
			end
			if(!(n7_odata_p0_21__gfpga === n7_odata_p0_21__bench) && !(n7_odata_p0_21__bench === 1'bx)) begin
				n7_odata_p0_21__flag <= 1'b1;
			end else begin
				n7_odata_p0_21__flag<= 1'b0;
			end
			if(!(n7_odata_p0_22__gfpga === n7_odata_p0_22__bench) && !(n7_odata_p0_22__bench === 1'bx)) begin
				n7_odata_p0_22__flag <= 1'b1;
			end else begin
				n7_odata_p0_22__flag<= 1'b0;
			end
			if(!(n7_odata_p0_23__gfpga === n7_odata_p0_23__bench) && !(n7_odata_p0_23__bench === 1'bx)) begin
				n7_odata_p0_23__flag <= 1'b1;
			end else begin
				n7_odata_p0_23__flag<= 1'b0;
			end
			if(!(n7_odata_p0_24__gfpga === n7_odata_p0_24__bench) && !(n7_odata_p0_24__bench === 1'bx)) begin
				n7_odata_p0_24__flag <= 1'b1;
			end else begin
				n7_odata_p0_24__flag<= 1'b0;
			end
			if(!(n7_odata_p0_25__gfpga === n7_odata_p0_25__bench) && !(n7_odata_p0_25__bench === 1'bx)) begin
				n7_odata_p0_25__flag <= 1'b1;
			end else begin
				n7_odata_p0_25__flag<= 1'b0;
			end
			if(!(n7_odata_p0_26__gfpga === n7_odata_p0_26__bench) && !(n7_odata_p0_26__bench === 1'bx)) begin
				n7_odata_p0_26__flag <= 1'b1;
			end else begin
				n7_odata_p0_26__flag<= 1'b0;
			end
			if(!(n7_odata_p0_27__gfpga === n7_odata_p0_27__bench) && !(n7_odata_p0_27__bench === 1'bx)) begin
				n7_odata_p0_27__flag <= 1'b1;
			end else begin
				n7_odata_p0_27__flag<= 1'b0;
			end
			if(!(n7_odata_p0_28__gfpga === n7_odata_p0_28__bench) && !(n7_odata_p0_28__bench === 1'bx)) begin
				n7_odata_p0_28__flag <= 1'b1;
			end else begin
				n7_odata_p0_28__flag<= 1'b0;
			end
			if(!(n7_odata_p0_29__gfpga === n7_odata_p0_29__bench) && !(n7_odata_p0_29__bench === 1'bx)) begin
				n7_odata_p0_29__flag <= 1'b1;
			end else begin
				n7_odata_p0_29__flag<= 1'b0;
			end
			if(!(n7_odata_p0_30__gfpga === n7_odata_p0_30__bench) && !(n7_odata_p0_30__bench === 1'bx)) begin
				n7_odata_p0_30__flag <= 1'b1;
			end else begin
				n7_odata_p0_30__flag<= 1'b0;
			end
			if(!(n7_odata_p0_31__gfpga === n7_odata_p0_31__bench) && !(n7_odata_p0_31__bench === 1'bx)) begin
				n7_odata_p0_31__flag <= 1'b1;
			end else begin
				n7_odata_p0_31__flag<= 1'b0;
			end
			if(!(n7_odata_p0_32__gfpga === n7_odata_p0_32__bench) && !(n7_odata_p0_32__bench === 1'bx)) begin
				n7_odata_p0_32__flag <= 1'b1;
			end else begin
				n7_odata_p0_32__flag<= 1'b0;
			end
			if(!(n7_odata_p0_33__gfpga === n7_odata_p0_33__bench) && !(n7_odata_p0_33__bench === 1'bx)) begin
				n7_odata_p0_33__flag <= 1'b1;
			end else begin
				n7_odata_p0_33__flag<= 1'b0;
			end
			if(!(n7_odata_p0_34__gfpga === n7_odata_p0_34__bench) && !(n7_odata_p0_34__bench === 1'bx)) begin
				n7_odata_p0_34__flag <= 1'b1;
			end else begin
				n7_odata_p0_34__flag<= 1'b0;
			end
			if(!(n7_ovalid_p0_gfpga === n7_ovalid_p0_bench) && !(n7_ovalid_p0_bench === 1'bx)) begin
				n7_ovalid_p0_flag <= 1'b1;
			end else begin
				n7_ovalid_p0_flag<= 1'b0;
			end
			if(!(n8_ordy_p0_0__gfpga === n8_ordy_p0_0__bench) && !(n8_ordy_p0_0__bench === 1'bx)) begin
				n8_ordy_p0_0__flag <= 1'b1;
			end else begin
				n8_ordy_p0_0__flag<= 1'b0;
			end
			if(!(n8_ordy_p0_1__gfpga === n8_ordy_p0_1__bench) && !(n8_ordy_p0_1__bench === 1'bx)) begin
				n8_ordy_p0_1__flag <= 1'b1;
			end else begin
				n8_ordy_p0_1__flag<= 1'b0;
			end
			if(!(n8_odata_p0_0__gfpga === n8_odata_p0_0__bench) && !(n8_odata_p0_0__bench === 1'bx)) begin
				n8_odata_p0_0__flag <= 1'b1;
			end else begin
				n8_odata_p0_0__flag<= 1'b0;
			end
			if(!(n8_odata_p0_1__gfpga === n8_odata_p0_1__bench) && !(n8_odata_p0_1__bench === 1'bx)) begin
				n8_odata_p0_1__flag <= 1'b1;
			end else begin
				n8_odata_p0_1__flag<= 1'b0;
			end
			if(!(n8_odata_p0_2__gfpga === n8_odata_p0_2__bench) && !(n8_odata_p0_2__bench === 1'bx)) begin
				n8_odata_p0_2__flag <= 1'b1;
			end else begin
				n8_odata_p0_2__flag<= 1'b0;
			end
			if(!(n8_odata_p0_3__gfpga === n8_odata_p0_3__bench) && !(n8_odata_p0_3__bench === 1'bx)) begin
				n8_odata_p0_3__flag <= 1'b1;
			end else begin
				n8_odata_p0_3__flag<= 1'b0;
			end
			if(!(n8_odata_p0_4__gfpga === n8_odata_p0_4__bench) && !(n8_odata_p0_4__bench === 1'bx)) begin
				n8_odata_p0_4__flag <= 1'b1;
			end else begin
				n8_odata_p0_4__flag<= 1'b0;
			end
			if(!(n8_odata_p0_5__gfpga === n8_odata_p0_5__bench) && !(n8_odata_p0_5__bench === 1'bx)) begin
				n8_odata_p0_5__flag <= 1'b1;
			end else begin
				n8_odata_p0_5__flag<= 1'b0;
			end
			if(!(n8_odata_p0_6__gfpga === n8_odata_p0_6__bench) && !(n8_odata_p0_6__bench === 1'bx)) begin
				n8_odata_p0_6__flag <= 1'b1;
			end else begin
				n8_odata_p0_6__flag<= 1'b0;
			end
			if(!(n8_odata_p0_7__gfpga === n8_odata_p0_7__bench) && !(n8_odata_p0_7__bench === 1'bx)) begin
				n8_odata_p0_7__flag <= 1'b1;
			end else begin
				n8_odata_p0_7__flag<= 1'b0;
			end
			if(!(n8_odata_p0_8__gfpga === n8_odata_p0_8__bench) && !(n8_odata_p0_8__bench === 1'bx)) begin
				n8_odata_p0_8__flag <= 1'b1;
			end else begin
				n8_odata_p0_8__flag<= 1'b0;
			end
			if(!(n8_odata_p0_9__gfpga === n8_odata_p0_9__bench) && !(n8_odata_p0_9__bench === 1'bx)) begin
				n8_odata_p0_9__flag <= 1'b1;
			end else begin
				n8_odata_p0_9__flag<= 1'b0;
			end
			if(!(n8_odata_p0_10__gfpga === n8_odata_p0_10__bench) && !(n8_odata_p0_10__bench === 1'bx)) begin
				n8_odata_p0_10__flag <= 1'b1;
			end else begin
				n8_odata_p0_10__flag<= 1'b0;
			end
			if(!(n8_odata_p0_11__gfpga === n8_odata_p0_11__bench) && !(n8_odata_p0_11__bench === 1'bx)) begin
				n8_odata_p0_11__flag <= 1'b1;
			end else begin
				n8_odata_p0_11__flag<= 1'b0;
			end
			if(!(n8_odata_p0_12__gfpga === n8_odata_p0_12__bench) && !(n8_odata_p0_12__bench === 1'bx)) begin
				n8_odata_p0_12__flag <= 1'b1;
			end else begin
				n8_odata_p0_12__flag<= 1'b0;
			end
			if(!(n8_odata_p0_13__gfpga === n8_odata_p0_13__bench) && !(n8_odata_p0_13__bench === 1'bx)) begin
				n8_odata_p0_13__flag <= 1'b1;
			end else begin
				n8_odata_p0_13__flag<= 1'b0;
			end
			if(!(n8_odata_p0_14__gfpga === n8_odata_p0_14__bench) && !(n8_odata_p0_14__bench === 1'bx)) begin
				n8_odata_p0_14__flag <= 1'b1;
			end else begin
				n8_odata_p0_14__flag<= 1'b0;
			end
			if(!(n8_odata_p0_15__gfpga === n8_odata_p0_15__bench) && !(n8_odata_p0_15__bench === 1'bx)) begin
				n8_odata_p0_15__flag <= 1'b1;
			end else begin
				n8_odata_p0_15__flag<= 1'b0;
			end
			if(!(n8_odata_p0_16__gfpga === n8_odata_p0_16__bench) && !(n8_odata_p0_16__bench === 1'bx)) begin
				n8_odata_p0_16__flag <= 1'b1;
			end else begin
				n8_odata_p0_16__flag<= 1'b0;
			end
			if(!(n8_odata_p0_17__gfpga === n8_odata_p0_17__bench) && !(n8_odata_p0_17__bench === 1'bx)) begin
				n8_odata_p0_17__flag <= 1'b1;
			end else begin
				n8_odata_p0_17__flag<= 1'b0;
			end
			if(!(n8_odata_p0_18__gfpga === n8_odata_p0_18__bench) && !(n8_odata_p0_18__bench === 1'bx)) begin
				n8_odata_p0_18__flag <= 1'b1;
			end else begin
				n8_odata_p0_18__flag<= 1'b0;
			end
			if(!(n8_odata_p0_19__gfpga === n8_odata_p0_19__bench) && !(n8_odata_p0_19__bench === 1'bx)) begin
				n8_odata_p0_19__flag <= 1'b1;
			end else begin
				n8_odata_p0_19__flag<= 1'b0;
			end
			if(!(n8_odata_p0_20__gfpga === n8_odata_p0_20__bench) && !(n8_odata_p0_20__bench === 1'bx)) begin
				n8_odata_p0_20__flag <= 1'b1;
			end else begin
				n8_odata_p0_20__flag<= 1'b0;
			end
			if(!(n8_odata_p0_21__gfpga === n8_odata_p0_21__bench) && !(n8_odata_p0_21__bench === 1'bx)) begin
				n8_odata_p0_21__flag <= 1'b1;
			end else begin
				n8_odata_p0_21__flag<= 1'b0;
			end
			if(!(n8_odata_p0_22__gfpga === n8_odata_p0_22__bench) && !(n8_odata_p0_22__bench === 1'bx)) begin
				n8_odata_p0_22__flag <= 1'b1;
			end else begin
				n8_odata_p0_22__flag<= 1'b0;
			end
			if(!(n8_odata_p0_23__gfpga === n8_odata_p0_23__bench) && !(n8_odata_p0_23__bench === 1'bx)) begin
				n8_odata_p0_23__flag <= 1'b1;
			end else begin
				n8_odata_p0_23__flag<= 1'b0;
			end
			if(!(n8_odata_p0_24__gfpga === n8_odata_p0_24__bench) && !(n8_odata_p0_24__bench === 1'bx)) begin
				n8_odata_p0_24__flag <= 1'b1;
			end else begin
				n8_odata_p0_24__flag<= 1'b0;
			end
			if(!(n8_odata_p0_25__gfpga === n8_odata_p0_25__bench) && !(n8_odata_p0_25__bench === 1'bx)) begin
				n8_odata_p0_25__flag <= 1'b1;
			end else begin
				n8_odata_p0_25__flag<= 1'b0;
			end
			if(!(n8_odata_p0_26__gfpga === n8_odata_p0_26__bench) && !(n8_odata_p0_26__bench === 1'bx)) begin
				n8_odata_p0_26__flag <= 1'b1;
			end else begin
				n8_odata_p0_26__flag<= 1'b0;
			end
			if(!(n8_odata_p0_27__gfpga === n8_odata_p0_27__bench) && !(n8_odata_p0_27__bench === 1'bx)) begin
				n8_odata_p0_27__flag <= 1'b1;
			end else begin
				n8_odata_p0_27__flag<= 1'b0;
			end
			if(!(n8_odata_p0_28__gfpga === n8_odata_p0_28__bench) && !(n8_odata_p0_28__bench === 1'bx)) begin
				n8_odata_p0_28__flag <= 1'b1;
			end else begin
				n8_odata_p0_28__flag<= 1'b0;
			end
			if(!(n8_odata_p0_29__gfpga === n8_odata_p0_29__bench) && !(n8_odata_p0_29__bench === 1'bx)) begin
				n8_odata_p0_29__flag <= 1'b1;
			end else begin
				n8_odata_p0_29__flag<= 1'b0;
			end
			if(!(n8_odata_p0_30__gfpga === n8_odata_p0_30__bench) && !(n8_odata_p0_30__bench === 1'bx)) begin
				n8_odata_p0_30__flag <= 1'b1;
			end else begin
				n8_odata_p0_30__flag<= 1'b0;
			end
			if(!(n8_odata_p0_31__gfpga === n8_odata_p0_31__bench) && !(n8_odata_p0_31__bench === 1'bx)) begin
				n8_odata_p0_31__flag <= 1'b1;
			end else begin
				n8_odata_p0_31__flag<= 1'b0;
			end
			if(!(n8_odata_p0_32__gfpga === n8_odata_p0_32__bench) && !(n8_odata_p0_32__bench === 1'bx)) begin
				n8_odata_p0_32__flag <= 1'b1;
			end else begin
				n8_odata_p0_32__flag<= 1'b0;
			end
			if(!(n8_odata_p0_33__gfpga === n8_odata_p0_33__bench) && !(n8_odata_p0_33__bench === 1'bx)) begin
				n8_odata_p0_33__flag <= 1'b1;
			end else begin
				n8_odata_p0_33__flag<= 1'b0;
			end
			if(!(n8_odata_p0_34__gfpga === n8_odata_p0_34__bench) && !(n8_odata_p0_34__bench === 1'bx)) begin
				n8_odata_p0_34__flag <= 1'b1;
			end else begin
				n8_odata_p0_34__flag<= 1'b0;
			end
			if(!(n8_ovalid_p0_gfpga === n8_ovalid_p0_bench) && !(n8_ovalid_p0_bench === 1'bx)) begin
				n8_ovalid_p0_flag <= 1'b1;
			end else begin
				n8_ovalid_p0_flag<= 1'b0;
			end
		end
	end

	always@(posedge n0_ordy_p0_0__flag) begin
		if(n0_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_ordy_p0_1__flag) begin
		if(n0_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_0__flag) begin
		if(n0_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_1__flag) begin
		if(n0_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_2__flag) begin
		if(n0_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_3__flag) begin
		if(n0_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_4__flag) begin
		if(n0_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_5__flag) begin
		if(n0_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_6__flag) begin
		if(n0_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_7__flag) begin
		if(n0_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_8__flag) begin
		if(n0_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_9__flag) begin
		if(n0_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_10__flag) begin
		if(n0_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_11__flag) begin
		if(n0_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_12__flag) begin
		if(n0_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_13__flag) begin
		if(n0_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_14__flag) begin
		if(n0_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_15__flag) begin
		if(n0_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_16__flag) begin
		if(n0_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_17__flag) begin
		if(n0_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_18__flag) begin
		if(n0_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_19__flag) begin
		if(n0_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_20__flag) begin
		if(n0_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_21__flag) begin
		if(n0_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_22__flag) begin
		if(n0_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_23__flag) begin
		if(n0_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_24__flag) begin
		if(n0_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_25__flag) begin
		if(n0_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_26__flag) begin
		if(n0_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_27__flag) begin
		if(n0_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_28__flag) begin
		if(n0_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_29__flag) begin
		if(n0_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_30__flag) begin
		if(n0_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_31__flag) begin
		if(n0_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_32__flag) begin
		if(n0_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_33__flag) begin
		if(n0_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_odata_p0_34__flag) begin
		if(n0_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n0_ovalid_p0_flag) begin
		if(n0_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n0_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_ordy_p0_0__flag) begin
		if(n1_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_ordy_p0_1__flag) begin
		if(n1_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_0__flag) begin
		if(n1_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_1__flag) begin
		if(n1_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_2__flag) begin
		if(n1_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_3__flag) begin
		if(n1_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_4__flag) begin
		if(n1_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_5__flag) begin
		if(n1_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_6__flag) begin
		if(n1_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_7__flag) begin
		if(n1_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_8__flag) begin
		if(n1_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_9__flag) begin
		if(n1_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_10__flag) begin
		if(n1_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_11__flag) begin
		if(n1_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_12__flag) begin
		if(n1_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_13__flag) begin
		if(n1_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_14__flag) begin
		if(n1_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_15__flag) begin
		if(n1_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_16__flag) begin
		if(n1_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_17__flag) begin
		if(n1_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_18__flag) begin
		if(n1_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_19__flag) begin
		if(n1_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_20__flag) begin
		if(n1_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_21__flag) begin
		if(n1_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_22__flag) begin
		if(n1_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_23__flag) begin
		if(n1_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_24__flag) begin
		if(n1_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_25__flag) begin
		if(n1_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_26__flag) begin
		if(n1_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_27__flag) begin
		if(n1_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_28__flag) begin
		if(n1_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_29__flag) begin
		if(n1_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_30__flag) begin
		if(n1_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_31__flag) begin
		if(n1_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_32__flag) begin
		if(n1_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_33__flag) begin
		if(n1_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_odata_p0_34__flag) begin
		if(n1_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n1_ovalid_p0_flag) begin
		if(n1_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n1_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_ordy_p0_0__flag) begin
		if(n2_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_ordy_p0_1__flag) begin
		if(n2_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_0__flag) begin
		if(n2_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_1__flag) begin
		if(n2_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_2__flag) begin
		if(n2_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_3__flag) begin
		if(n2_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_4__flag) begin
		if(n2_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_5__flag) begin
		if(n2_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_6__flag) begin
		if(n2_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_7__flag) begin
		if(n2_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_8__flag) begin
		if(n2_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_9__flag) begin
		if(n2_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_10__flag) begin
		if(n2_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_11__flag) begin
		if(n2_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_12__flag) begin
		if(n2_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_13__flag) begin
		if(n2_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_14__flag) begin
		if(n2_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_15__flag) begin
		if(n2_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_16__flag) begin
		if(n2_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_17__flag) begin
		if(n2_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_18__flag) begin
		if(n2_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_19__flag) begin
		if(n2_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_20__flag) begin
		if(n2_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_21__flag) begin
		if(n2_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_22__flag) begin
		if(n2_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_23__flag) begin
		if(n2_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_24__flag) begin
		if(n2_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_25__flag) begin
		if(n2_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_26__flag) begin
		if(n2_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_27__flag) begin
		if(n2_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_28__flag) begin
		if(n2_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_29__flag) begin
		if(n2_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_30__flag) begin
		if(n2_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_31__flag) begin
		if(n2_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_32__flag) begin
		if(n2_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_33__flag) begin
		if(n2_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_odata_p0_34__flag) begin
		if(n2_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n2_ovalid_p0_flag) begin
		if(n2_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n2_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_ordy_p0_0__flag) begin
		if(n3_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_ordy_p0_1__flag) begin
		if(n3_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_0__flag) begin
		if(n3_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_1__flag) begin
		if(n3_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_2__flag) begin
		if(n3_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_3__flag) begin
		if(n3_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_4__flag) begin
		if(n3_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_5__flag) begin
		if(n3_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_6__flag) begin
		if(n3_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_7__flag) begin
		if(n3_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_8__flag) begin
		if(n3_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_9__flag) begin
		if(n3_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_10__flag) begin
		if(n3_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_11__flag) begin
		if(n3_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_12__flag) begin
		if(n3_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_13__flag) begin
		if(n3_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_14__flag) begin
		if(n3_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_15__flag) begin
		if(n3_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_16__flag) begin
		if(n3_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_17__flag) begin
		if(n3_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_18__flag) begin
		if(n3_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_19__flag) begin
		if(n3_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_20__flag) begin
		if(n3_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_21__flag) begin
		if(n3_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_22__flag) begin
		if(n3_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_23__flag) begin
		if(n3_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_24__flag) begin
		if(n3_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_25__flag) begin
		if(n3_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_26__flag) begin
		if(n3_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_27__flag) begin
		if(n3_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_28__flag) begin
		if(n3_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_29__flag) begin
		if(n3_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_30__flag) begin
		if(n3_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_31__flag) begin
		if(n3_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_32__flag) begin
		if(n3_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_33__flag) begin
		if(n3_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_odata_p0_34__flag) begin
		if(n3_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n3_ovalid_p0_flag) begin
		if(n3_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n3_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_ordy_p0_0__flag) begin
		if(n4_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_ordy_p0_1__flag) begin
		if(n4_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_0__flag) begin
		if(n4_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_1__flag) begin
		if(n4_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_2__flag) begin
		if(n4_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_3__flag) begin
		if(n4_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_4__flag) begin
		if(n4_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_5__flag) begin
		if(n4_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_6__flag) begin
		if(n4_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_7__flag) begin
		if(n4_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_8__flag) begin
		if(n4_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_9__flag) begin
		if(n4_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_10__flag) begin
		if(n4_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_11__flag) begin
		if(n4_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_12__flag) begin
		if(n4_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_13__flag) begin
		if(n4_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_14__flag) begin
		if(n4_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_15__flag) begin
		if(n4_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_16__flag) begin
		if(n4_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_17__flag) begin
		if(n4_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_18__flag) begin
		if(n4_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_19__flag) begin
		if(n4_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_20__flag) begin
		if(n4_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_21__flag) begin
		if(n4_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_22__flag) begin
		if(n4_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_23__flag) begin
		if(n4_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_24__flag) begin
		if(n4_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_25__flag) begin
		if(n4_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_26__flag) begin
		if(n4_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_27__flag) begin
		if(n4_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_28__flag) begin
		if(n4_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_29__flag) begin
		if(n4_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_30__flag) begin
		if(n4_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_31__flag) begin
		if(n4_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_32__flag) begin
		if(n4_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_33__flag) begin
		if(n4_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_odata_p0_34__flag) begin
		if(n4_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n4_ovalid_p0_flag) begin
		if(n4_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n4_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_ordy_p0_0__flag) begin
		if(n5_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_ordy_p0_1__flag) begin
		if(n5_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_0__flag) begin
		if(n5_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_1__flag) begin
		if(n5_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_2__flag) begin
		if(n5_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_3__flag) begin
		if(n5_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_4__flag) begin
		if(n5_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_5__flag) begin
		if(n5_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_6__flag) begin
		if(n5_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_7__flag) begin
		if(n5_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_8__flag) begin
		if(n5_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_9__flag) begin
		if(n5_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_10__flag) begin
		if(n5_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_11__flag) begin
		if(n5_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_12__flag) begin
		if(n5_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_13__flag) begin
		if(n5_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_14__flag) begin
		if(n5_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_15__flag) begin
		if(n5_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_16__flag) begin
		if(n5_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_17__flag) begin
		if(n5_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_18__flag) begin
		if(n5_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_19__flag) begin
		if(n5_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_20__flag) begin
		if(n5_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_21__flag) begin
		if(n5_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_22__flag) begin
		if(n5_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_23__flag) begin
		if(n5_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_24__flag) begin
		if(n5_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_25__flag) begin
		if(n5_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_26__flag) begin
		if(n5_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_27__flag) begin
		if(n5_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_28__flag) begin
		if(n5_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_29__flag) begin
		if(n5_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_30__flag) begin
		if(n5_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_31__flag) begin
		if(n5_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_32__flag) begin
		if(n5_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_33__flag) begin
		if(n5_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_odata_p0_34__flag) begin
		if(n5_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n5_ovalid_p0_flag) begin
		if(n5_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n5_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_ordy_p0_0__flag) begin
		if(n6_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_ordy_p0_1__flag) begin
		if(n6_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_0__flag) begin
		if(n6_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_1__flag) begin
		if(n6_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_2__flag) begin
		if(n6_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_3__flag) begin
		if(n6_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_4__flag) begin
		if(n6_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_5__flag) begin
		if(n6_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_6__flag) begin
		if(n6_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_7__flag) begin
		if(n6_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_8__flag) begin
		if(n6_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_9__flag) begin
		if(n6_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_10__flag) begin
		if(n6_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_11__flag) begin
		if(n6_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_12__flag) begin
		if(n6_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_13__flag) begin
		if(n6_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_14__flag) begin
		if(n6_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_15__flag) begin
		if(n6_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_16__flag) begin
		if(n6_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_17__flag) begin
		if(n6_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_18__flag) begin
		if(n6_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_19__flag) begin
		if(n6_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_20__flag) begin
		if(n6_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_21__flag) begin
		if(n6_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_22__flag) begin
		if(n6_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_23__flag) begin
		if(n6_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_24__flag) begin
		if(n6_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_25__flag) begin
		if(n6_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_26__flag) begin
		if(n6_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_27__flag) begin
		if(n6_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_28__flag) begin
		if(n6_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_29__flag) begin
		if(n6_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_30__flag) begin
		if(n6_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_31__flag) begin
		if(n6_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_32__flag) begin
		if(n6_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_33__flag) begin
		if(n6_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_odata_p0_34__flag) begin
		if(n6_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n6_ovalid_p0_flag) begin
		if(n6_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n6_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_ordy_p0_0__flag) begin
		if(n7_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_ordy_p0_1__flag) begin
		if(n7_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_0__flag) begin
		if(n7_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_1__flag) begin
		if(n7_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_2__flag) begin
		if(n7_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_3__flag) begin
		if(n7_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_4__flag) begin
		if(n7_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_5__flag) begin
		if(n7_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_6__flag) begin
		if(n7_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_7__flag) begin
		if(n7_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_8__flag) begin
		if(n7_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_9__flag) begin
		if(n7_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_10__flag) begin
		if(n7_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_11__flag) begin
		if(n7_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_12__flag) begin
		if(n7_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_13__flag) begin
		if(n7_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_14__flag) begin
		if(n7_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_15__flag) begin
		if(n7_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_16__flag) begin
		if(n7_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_17__flag) begin
		if(n7_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_18__flag) begin
		if(n7_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_19__flag) begin
		if(n7_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_20__flag) begin
		if(n7_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_21__flag) begin
		if(n7_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_22__flag) begin
		if(n7_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_23__flag) begin
		if(n7_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_24__flag) begin
		if(n7_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_25__flag) begin
		if(n7_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_26__flag) begin
		if(n7_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_27__flag) begin
		if(n7_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_28__flag) begin
		if(n7_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_29__flag) begin
		if(n7_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_30__flag) begin
		if(n7_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_31__flag) begin
		if(n7_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_32__flag) begin
		if(n7_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_33__flag) begin
		if(n7_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_odata_p0_34__flag) begin
		if(n7_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n7_ovalid_p0_flag) begin
		if(n7_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n7_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_ordy_p0_0__flag) begin
		if(n8_ordy_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_ordy_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_ordy_p0_1__flag) begin
		if(n8_ordy_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_ordy_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_0__flag) begin
		if(n8_odata_p0_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_1__flag) begin
		if(n8_odata_p0_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_2__flag) begin
		if(n8_odata_p0_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_3__flag) begin
		if(n8_odata_p0_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_4__flag) begin
		if(n8_odata_p0_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_5__flag) begin
		if(n8_odata_p0_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_6__flag) begin
		if(n8_odata_p0_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_7__flag) begin
		if(n8_odata_p0_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_8__flag) begin
		if(n8_odata_p0_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_9__flag) begin
		if(n8_odata_p0_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_10__flag) begin
		if(n8_odata_p0_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_11__flag) begin
		if(n8_odata_p0_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_12__flag) begin
		if(n8_odata_p0_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_13__flag) begin
		if(n8_odata_p0_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_14__flag) begin
		if(n8_odata_p0_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_15__flag) begin
		if(n8_odata_p0_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_16__flag) begin
		if(n8_odata_p0_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_17__flag) begin
		if(n8_odata_p0_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_18__flag) begin
		if(n8_odata_p0_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_19__flag) begin
		if(n8_odata_p0_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_20__flag) begin
		if(n8_odata_p0_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_21__flag) begin
		if(n8_odata_p0_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_22__flag) begin
		if(n8_odata_p0_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_23__flag) begin
		if(n8_odata_p0_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_24__flag) begin
		if(n8_odata_p0_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_25__flag) begin
		if(n8_odata_p0_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_26__flag) begin
		if(n8_odata_p0_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_27__flag) begin
		if(n8_odata_p0_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_28__flag) begin
		if(n8_odata_p0_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_29__flag) begin
		if(n8_odata_p0_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_30__flag) begin
		if(n8_odata_p0_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_31__flag) begin
		if(n8_odata_p0_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_32__flag) begin
		if(n8_odata_p0_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_33__flag) begin
		if(n8_odata_p0_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_odata_p0_34__flag) begin
		if(n8_odata_p0_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_odata_p0_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge n8_ovalid_p0_flag) begin
		if(n8_ovalid_p0_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on n8_ovalid_p0_gfpga at time = %t", $realtime);
		end
	end


// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("noc_formal.vcd");
		$dumpvars(1, noc_top_formal_verification_random_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#20
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for noc_top_formal_verification_random_tb -----

