//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: mesh_bench
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Aug  8 17:59:29 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module mesh_bench_top_formal_verification (
input [0:0] i_data_0_0_,
input [0:0] i_data_0_1_,
input [0:0] i_data_0_2_,
input [0:0] i_data_0_3_,
input [0:0] i_data_0_4_,
input [0:0] i_data_0_5_,
input [0:0] i_data_0_6_,
input [0:0] i_data_0_7_,
input [0:0] i_data_0_8_,
input [0:0] i_data_0_9_,
input [0:0] i_data_0_10_,
input [0:0] i_data_0_11_,
input [0:0] i_data_0_12_,
input [0:0] i_data_0_13_,
input [0:0] i_data_0_14_,
input [0:0] i_data_0_15_,
input [0:0] i_data_0_16_,
input [0:0] i_data_0_17_,
input [0:0] i_data_0_18_,
input [0:0] i_data_0_19_,
input [0:0] i_data_0_20_,
input [0:0] i_data_0_21_,
input [0:0] i_data_0_22_,
input [0:0] i_data_0_23_,
input [0:0] i_data_0_24_,
input [0:0] i_data_0_25_,
input [0:0] i_data_0_26_,
input [0:0] i_data_0_27_,
input [0:0] i_data_0_28_,
input [0:0] i_data_0_29_,
input [0:0] i_data_0_30_,
input [0:0] i_data_0_31_,
input [0:0] i_data_0_32_,
input [0:0] i_data_0_33_,
input [0:0] i_data_0_34_,
input [0:0] i_valid_0,
input [0:0] i_vch_0,
input [0:0] i_ack_0_0_,
input [0:0] i_ack_0_1_,
input [0:0] i_lck_0_0_,
input [0:0] i_lck_0_1_,
input [0:0] i_data_1_0_,
input [0:0] i_data_1_1_,
input [0:0] i_data_1_2_,
input [0:0] i_data_1_3_,
input [0:0] i_data_1_4_,
input [0:0] i_data_1_5_,
input [0:0] i_data_1_6_,
input [0:0] i_data_1_7_,
input [0:0] i_data_1_8_,
input [0:0] i_data_1_9_,
input [0:0] i_data_1_10_,
input [0:0] i_data_1_11_,
input [0:0] i_data_1_12_,
input [0:0] i_data_1_13_,
input [0:0] i_data_1_14_,
input [0:0] i_data_1_15_,
input [0:0] i_data_1_16_,
input [0:0] i_data_1_17_,
input [0:0] i_data_1_18_,
input [0:0] i_data_1_19_,
input [0:0] i_data_1_20_,
input [0:0] i_data_1_21_,
input [0:0] i_data_1_22_,
input [0:0] i_data_1_23_,
input [0:0] i_data_1_24_,
input [0:0] i_data_1_25_,
input [0:0] i_data_1_26_,
input [0:0] i_data_1_27_,
input [0:0] i_data_1_28_,
input [0:0] i_data_1_29_,
input [0:0] i_data_1_30_,
input [0:0] i_data_1_31_,
input [0:0] i_data_1_32_,
input [0:0] i_data_1_33_,
input [0:0] i_data_1_34_,
input [0:0] i_valid_1,
input [0:0] i_vch_1,
input [0:0] i_ack_1_0_,
input [0:0] i_ack_1_1_,
input [0:0] i_lck_1_0_,
input [0:0] i_lck_1_1_,
input [0:0] clk,
input [0:0] rst_,
output [0:0] o_data_0_0_,
output [0:0] o_data_0_1_,
output [0:0] o_data_0_2_,
output [0:0] o_data_0_3_,
output [0:0] o_data_0_4_,
output [0:0] o_data_0_5_,
output [0:0] o_data_0_6_,
output [0:0] o_data_0_7_,
output [0:0] o_data_0_8_,
output [0:0] o_data_0_9_,
output [0:0] o_data_0_10_,
output [0:0] o_data_0_11_,
output [0:0] o_data_0_12_,
output [0:0] o_data_0_13_,
output [0:0] o_data_0_14_,
output [0:0] o_data_0_15_,
output [0:0] o_data_0_16_,
output [0:0] o_data_0_17_,
output [0:0] o_data_0_18_,
output [0:0] o_data_0_19_,
output [0:0] o_data_0_20_,
output [0:0] o_data_0_21_,
output [0:0] o_data_0_22_,
output [0:0] o_data_0_23_,
output [0:0] o_data_0_24_,
output [0:0] o_data_0_25_,
output [0:0] o_data_0_26_,
output [0:0] o_data_0_27_,
output [0:0] o_data_0_28_,
output [0:0] o_data_0_29_,
output [0:0] o_data_0_30_,
output [0:0] o_data_0_31_,
output [0:0] o_data_0_32_,
output [0:0] o_data_0_33_,
output [0:0] o_data_0_34_,
output [0:0] o_valid_0,
output [0:0] o_vch_0,
output [0:0] o_ack_0_0_,
output [0:0] o_ack_0_1_,
output [0:0] o_lck_0_0_,
output [0:0] o_lck_0_1_,
output [0:0] o_rdy_0_0_,
output [0:0] o_rdy_0_1_,
output [0:0] o_data_1_0_,
output [0:0] o_data_1_1_,
output [0:0] o_data_1_2_,
output [0:0] o_data_1_3_,
output [0:0] o_data_1_4_,
output [0:0] o_data_1_5_,
output [0:0] o_data_1_6_,
output [0:0] o_data_1_7_,
output [0:0] o_data_1_8_,
output [0:0] o_data_1_9_,
output [0:0] o_data_1_10_,
output [0:0] o_data_1_11_,
output [0:0] o_data_1_12_,
output [0:0] o_data_1_13_,
output [0:0] o_data_1_14_,
output [0:0] o_data_1_15_,
output [0:0] o_data_1_16_,
output [0:0] o_data_1_17_,
output [0:0] o_data_1_18_,
output [0:0] o_data_1_19_,
output [0:0] o_data_1_20_,
output [0:0] o_data_1_21_,
output [0:0] o_data_1_22_,
output [0:0] o_data_1_23_,
output [0:0] o_data_1_24_,
output [0:0] o_data_1_25_,
output [0:0] o_data_1_26_,
output [0:0] o_data_1_27_,
output [0:0] o_data_1_28_,
output [0:0] o_data_1_29_,
output [0:0] o_data_1_30_,
output [0:0] o_data_1_31_,
output [0:0] o_data_1_32_,
output [0:0] o_data_1_33_,
output [0:0] o_data_1_34_,
output [0:0] o_valid_1,
output [0:0] o_vch_1,
output [0:0] o_ack_1_0_,
output [0:0] o_ack_1_1_,
output [0:0] o_lck_1_0_,
output [0:0] o_lck_1_1_,
output [0:0] o_rdy_1_0_,
output [0:0] o_rdy_1_1_);

// ----- Local wires for FPGA fabric -----
wire [0:223] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] pReset_fm;
wire [0:0] prog_clk_fm;
wire [0:0] clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		pReset_fm[0],
		prog_clk_fm[0],
		clk_fm[0],
		set_fm[0],
		reset_fm[0],
		gfpga_pad_GPIO_PAD_fm[0:223],
		ccff_head_fm[0],
		ccff_tail_fm[0]);

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = 1'b0;
	assign clk_fm[0] = clk[0];
	assign pReset_fm[0] = 1'b0;
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input i_data_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[103] -----
	assign gfpga_pad_GPIO_PAD_fm[103] = i_data_0_0_[0];

// ----- Blif Benchmark input i_data_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[102] -----
	assign gfpga_pad_GPIO_PAD_fm[102] = i_data_0_1_[0];

// ----- Blif Benchmark input i_data_0_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[93] -----
	assign gfpga_pad_GPIO_PAD_fm[93] = i_data_0_2_[0];

// ----- Blif Benchmark input i_data_0_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[124] -----
	assign gfpga_pad_GPIO_PAD_fm[124] = i_data_0_3_[0];

// ----- Blif Benchmark input i_data_0_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[65] -----
	assign gfpga_pad_GPIO_PAD_fm[65] = i_data_0_4_[0];

// ----- Blif Benchmark input i_data_0_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[66] -----
	assign gfpga_pad_GPIO_PAD_fm[66] = i_data_0_5_[0];

// ----- Blif Benchmark input i_data_0_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[146] -----
	assign gfpga_pad_GPIO_PAD_fm[146] = i_data_0_6_[0];

// ----- Blif Benchmark input i_data_0_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[73] -----
	assign gfpga_pad_GPIO_PAD_fm[73] = i_data_0_7_[0];

// ----- Blif Benchmark input i_data_0_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[125] -----
	assign gfpga_pad_GPIO_PAD_fm[125] = i_data_0_8_[0];

// ----- Blif Benchmark input i_data_0_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[56] -----
	assign gfpga_pad_GPIO_PAD_fm[56] = i_data_0_9_[0];

// ----- Blif Benchmark input i_data_0_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[130] -----
	assign gfpga_pad_GPIO_PAD_fm[130] = i_data_0_10_[0];

// ----- Blif Benchmark input i_data_0_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[77] -----
	assign gfpga_pad_GPIO_PAD_fm[77] = i_data_0_11_[0];

// ----- Blif Benchmark input i_data_0_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[112] -----
	assign gfpga_pad_GPIO_PAD_fm[112] = i_data_0_12_[0];

// ----- Blif Benchmark input i_data_0_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[74] -----
	assign gfpga_pad_GPIO_PAD_fm[74] = i_data_0_13_[0];

// ----- Blif Benchmark input i_data_0_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[140] -----
	assign gfpga_pad_GPIO_PAD_fm[140] = i_data_0_14_[0];

// ----- Blif Benchmark input i_data_0_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[133] -----
	assign gfpga_pad_GPIO_PAD_fm[133] = i_data_0_15_[0];

// ----- Blif Benchmark input i_data_0_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[106] -----
	assign gfpga_pad_GPIO_PAD_fm[106] = i_data_0_16_[0];

// ----- Blif Benchmark input i_data_0_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[86] -----
	assign gfpga_pad_GPIO_PAD_fm[86] = i_data_0_17_[0];

// ----- Blif Benchmark input i_data_0_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[135] -----
	assign gfpga_pad_GPIO_PAD_fm[135] = i_data_0_18_[0];

// ----- Blif Benchmark input i_data_0_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[75] -----
	assign gfpga_pad_GPIO_PAD_fm[75] = i_data_0_19_[0];

// ----- Blif Benchmark input i_data_0_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[128] -----
	assign gfpga_pad_GPIO_PAD_fm[128] = i_data_0_20_[0];

// ----- Blif Benchmark input i_data_0_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[118] -----
	assign gfpga_pad_GPIO_PAD_fm[118] = i_data_0_21_[0];

// ----- Blif Benchmark input i_data_0_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[80] -----
	assign gfpga_pad_GPIO_PAD_fm[80] = i_data_0_22_[0];

// ----- Blif Benchmark input i_data_0_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[116] -----
	assign gfpga_pad_GPIO_PAD_fm[116] = i_data_0_23_[0];

// ----- Blif Benchmark input i_data_0_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[114] -----
	assign gfpga_pad_GPIO_PAD_fm[114] = i_data_0_24_[0];

// ----- Blif Benchmark input i_data_0_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[95] -----
	assign gfpga_pad_GPIO_PAD_fm[95] = i_data_0_25_[0];

// ----- Blif Benchmark input i_data_0_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[76] -----
	assign gfpga_pad_GPIO_PAD_fm[76] = i_data_0_26_[0];

// ----- Blif Benchmark input i_data_0_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[71] -----
	assign gfpga_pad_GPIO_PAD_fm[71] = i_data_0_27_[0];

// ----- Blif Benchmark input i_data_0_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[129] -----
	assign gfpga_pad_GPIO_PAD_fm[129] = i_data_0_28_[0];

// ----- Blif Benchmark input i_data_0_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[105] -----
	assign gfpga_pad_GPIO_PAD_fm[105] = i_data_0_29_[0];

// ----- Blif Benchmark input i_data_0_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[107] -----
	assign gfpga_pad_GPIO_PAD_fm[107] = i_data_0_30_[0];

// ----- Blif Benchmark input i_data_0_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[141] -----
	assign gfpga_pad_GPIO_PAD_fm[141] = i_data_0_31_[0];

// ----- Blif Benchmark input i_data_0_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[62] -----
	assign gfpga_pad_GPIO_PAD_fm[62] = i_data_0_32_[0];

// ----- Blif Benchmark input i_data_0_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[121] -----
	assign gfpga_pad_GPIO_PAD_fm[121] = i_data_0_33_[0];

// ----- Blif Benchmark input i_data_0_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[98] -----
	assign gfpga_pad_GPIO_PAD_fm[98] = i_data_0_34_[0];

// ----- Blif Benchmark input i_valid_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[72] -----
	assign gfpga_pad_GPIO_PAD_fm[72] = i_valid_0[0];

// ----- Blif Benchmark input i_vch_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[131] -----
	assign gfpga_pad_GPIO_PAD_fm[131] = i_vch_0[0];

// ----- Blif Benchmark input i_ack_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[126] -----
	assign gfpga_pad_GPIO_PAD_fm[126] = i_ack_0_0_[0];

// ----- Blif Benchmark input i_ack_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[139] -----
	assign gfpga_pad_GPIO_PAD_fm[139] = i_ack_0_1_[0];

// ----- Blif Benchmark input i_lck_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[115] -----
	assign gfpga_pad_GPIO_PAD_fm[115] = i_lck_0_0_[0];

// ----- Blif Benchmark input i_lck_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[104] -----
	assign gfpga_pad_GPIO_PAD_fm[104] = i_lck_0_1_[0];

// ----- Blif Benchmark input i_data_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[221] -----
	assign gfpga_pad_GPIO_PAD_fm[221] = i_data_1_0_[0];

// ----- Blif Benchmark input i_data_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[210] -----
	assign gfpga_pad_GPIO_PAD_fm[210] = i_data_1_1_[0];

// ----- Blif Benchmark input i_data_1_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[192] -----
	assign gfpga_pad_GPIO_PAD_fm[192] = i_data_1_2_[0];

// ----- Blif Benchmark input i_data_1_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[4] -----
	assign gfpga_pad_GPIO_PAD_fm[4] = i_data_1_3_[0];

// ----- Blif Benchmark input i_data_1_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[199] -----
	assign gfpga_pad_GPIO_PAD_fm[199] = i_data_1_4_[0];

// ----- Blif Benchmark input i_data_1_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[19] -----
	assign gfpga_pad_GPIO_PAD_fm[19] = i_data_1_5_[0];

// ----- Blif Benchmark input i_data_1_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[204] -----
	assign gfpga_pad_GPIO_PAD_fm[204] = i_data_1_6_[0];

// ----- Blif Benchmark input i_data_1_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[3] -----
	assign gfpga_pad_GPIO_PAD_fm[3] = i_data_1_7_[0];

// ----- Blif Benchmark input i_data_1_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[203] -----
	assign gfpga_pad_GPIO_PAD_fm[203] = i_data_1_8_[0];

// ----- Blif Benchmark input i_data_1_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[194] -----
	assign gfpga_pad_GPIO_PAD_fm[194] = i_data_1_9_[0];

// ----- Blif Benchmark input i_data_1_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[163] -----
	assign gfpga_pad_GPIO_PAD_fm[163] = i_data_1_10_[0];

// ----- Blif Benchmark input i_data_1_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[193] -----
	assign gfpga_pad_GPIO_PAD_fm[193] = i_data_1_11_[0];

// ----- Blif Benchmark input i_data_1_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[2] -----
	assign gfpga_pad_GPIO_PAD_fm[2] = i_data_1_12_[0];

// ----- Blif Benchmark input i_data_1_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[198] -----
	assign gfpga_pad_GPIO_PAD_fm[198] = i_data_1_13_[0];

// ----- Blif Benchmark input i_data_1_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[196] -----
	assign gfpga_pad_GPIO_PAD_fm[196] = i_data_1_14_[0];

// ----- Blif Benchmark input i_data_1_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[213] -----
	assign gfpga_pad_GPIO_PAD_fm[213] = i_data_1_15_[0];

// ----- Blif Benchmark input i_data_1_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[215] -----
	assign gfpga_pad_GPIO_PAD_fm[215] = i_data_1_16_[0];

// ----- Blif Benchmark input i_data_1_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[216] -----
	assign gfpga_pad_GPIO_PAD_fm[216] = i_data_1_17_[0];

// ----- Blif Benchmark input i_data_1_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[205] -----
	assign gfpga_pad_GPIO_PAD_fm[205] = i_data_1_18_[0];

// ----- Blif Benchmark input i_data_1_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[201] -----
	assign gfpga_pad_GPIO_PAD_fm[201] = i_data_1_19_[0];

// ----- Blif Benchmark input i_data_1_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[208] -----
	assign gfpga_pad_GPIO_PAD_fm[208] = i_data_1_20_[0];

// ----- Blif Benchmark input i_data_1_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[207] -----
	assign gfpga_pad_GPIO_PAD_fm[207] = i_data_1_21_[0];

// ----- Blif Benchmark input i_data_1_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[223] -----
	assign gfpga_pad_GPIO_PAD_fm[223] = i_data_1_22_[0];

// ----- Blif Benchmark input i_data_1_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[200] -----
	assign gfpga_pad_GPIO_PAD_fm[200] = i_data_1_23_[0];

// ----- Blif Benchmark input i_data_1_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[218] -----
	assign gfpga_pad_GPIO_PAD_fm[218] = i_data_1_24_[0];

// ----- Blif Benchmark input i_data_1_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[206] -----
	assign gfpga_pad_GPIO_PAD_fm[206] = i_data_1_25_[0];

// ----- Blif Benchmark input i_data_1_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[7] -----
	assign gfpga_pad_GPIO_PAD_fm[7] = i_data_1_26_[0];

// ----- Blif Benchmark input i_data_1_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[160] -----
	assign gfpga_pad_GPIO_PAD_fm[160] = i_data_1_27_[0];

// ----- Blif Benchmark input i_data_1_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[6] -----
	assign gfpga_pad_GPIO_PAD_fm[6] = i_data_1_28_[0];

// ----- Blif Benchmark input i_data_1_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[212] -----
	assign gfpga_pad_GPIO_PAD_fm[212] = i_data_1_29_[0];

// ----- Blif Benchmark input i_data_1_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[161] -----
	assign gfpga_pad_GPIO_PAD_fm[161] = i_data_1_30_[0];

// ----- Blif Benchmark input i_data_1_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[202] -----
	assign gfpga_pad_GPIO_PAD_fm[202] = i_data_1_31_[0];

// ----- Blif Benchmark input i_data_1_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[217] -----
	assign gfpga_pad_GPIO_PAD_fm[217] = i_data_1_32_[0];

// ----- Blif Benchmark input i_data_1_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[219] -----
	assign gfpga_pad_GPIO_PAD_fm[219] = i_data_1_33_[0];

// ----- Blif Benchmark input i_data_1_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[220] -----
	assign gfpga_pad_GPIO_PAD_fm[220] = i_data_1_34_[0];

// ----- Blif Benchmark input i_valid_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[209] -----
	assign gfpga_pad_GPIO_PAD_fm[209] = i_valid_1[0];

// ----- Blif Benchmark input i_vch_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[211] -----
	assign gfpga_pad_GPIO_PAD_fm[211] = i_vch_1[0];

// ----- Blif Benchmark input i_ack_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[195] -----
	assign gfpga_pad_GPIO_PAD_fm[195] = i_ack_1_0_[0];

// ----- Blif Benchmark input i_ack_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[214] -----
	assign gfpga_pad_GPIO_PAD_fm[214] = i_ack_1_1_[0];

// ----- Blif Benchmark input i_lck_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[222] -----
	assign gfpga_pad_GPIO_PAD_fm[222] = i_lck_1_0_[0];

// ----- Blif Benchmark input i_lck_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[167] -----
	assign gfpga_pad_GPIO_PAD_fm[167] = i_lck_1_1_[0];

// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[14] -----
	assign gfpga_pad_GPIO_PAD_fm[14] = clk[0];

// ----- Blif Benchmark input rst_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[151] -----
	assign gfpga_pad_GPIO_PAD_fm[151] = rst_[0];

// ----- Blif Benchmark output o_data_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[113] -----
	assign o_data_0_0_[0] = gfpga_pad_GPIO_PAD_fm[113];

// ----- Blif Benchmark output o_data_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[111] -----
	assign o_data_0_1_[0] = gfpga_pad_GPIO_PAD_fm[111];

// ----- Blif Benchmark output o_data_0_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[136] -----
	assign o_data_0_2_[0] = gfpga_pad_GPIO_PAD_fm[136];

// ----- Blif Benchmark output o_data_0_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[68] -----
	assign o_data_0_3_[0] = gfpga_pad_GPIO_PAD_fm[68];

// ----- Blif Benchmark output o_data_0_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[79] -----
	assign o_data_0_4_[0] = gfpga_pad_GPIO_PAD_fm[79];

// ----- Blif Benchmark output o_data_0_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[122] -----
	assign o_data_0_5_[0] = gfpga_pad_GPIO_PAD_fm[122];

// ----- Blif Benchmark output o_data_0_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[89] -----
	assign o_data_0_6_[0] = gfpga_pad_GPIO_PAD_fm[89];

// ----- Blif Benchmark output o_data_0_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[94] -----
	assign o_data_0_7_[0] = gfpga_pad_GPIO_PAD_fm[94];

// ----- Blif Benchmark output o_data_0_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[134] -----
	assign o_data_0_8_[0] = gfpga_pad_GPIO_PAD_fm[134];

// ----- Blif Benchmark output o_data_0_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[109] -----
	assign o_data_0_9_[0] = gfpga_pad_GPIO_PAD_fm[109];

// ----- Blif Benchmark output o_data_0_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[96] -----
	assign o_data_0_10_[0] = gfpga_pad_GPIO_PAD_fm[96];

// ----- Blif Benchmark output o_data_0_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[84] -----
	assign o_data_0_11_[0] = gfpga_pad_GPIO_PAD_fm[84];

// ----- Blif Benchmark output o_data_0_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[91] -----
	assign o_data_0_12_[0] = gfpga_pad_GPIO_PAD_fm[91];

// ----- Blif Benchmark output o_data_0_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[88] -----
	assign o_data_0_13_[0] = gfpga_pad_GPIO_PAD_fm[88];

// ----- Blif Benchmark output o_data_0_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[99] -----
	assign o_data_0_14_[0] = gfpga_pad_GPIO_PAD_fm[99];

// ----- Blif Benchmark output o_data_0_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[78] -----
	assign o_data_0_15_[0] = gfpga_pad_GPIO_PAD_fm[78];

// ----- Blif Benchmark output o_data_0_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[123] -----
	assign o_data_0_16_[0] = gfpga_pad_GPIO_PAD_fm[123];

// ----- Blif Benchmark output o_data_0_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[67] -----
	assign o_data_0_17_[0] = gfpga_pad_GPIO_PAD_fm[67];

// ----- Blif Benchmark output o_data_0_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[70] -----
	assign o_data_0_18_[0] = gfpga_pad_GPIO_PAD_fm[70];

// ----- Blif Benchmark output o_data_0_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[138] -----
	assign o_data_0_19_[0] = gfpga_pad_GPIO_PAD_fm[138];

// ----- Blif Benchmark output o_data_0_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[87] -----
	assign o_data_0_20_[0] = gfpga_pad_GPIO_PAD_fm[87];

// ----- Blif Benchmark output o_data_0_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[85] -----
	assign o_data_0_21_[0] = gfpga_pad_GPIO_PAD_fm[85];

// ----- Blif Benchmark output o_data_0_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[81] -----
	assign o_data_0_22_[0] = gfpga_pad_GPIO_PAD_fm[81];

// ----- Blif Benchmark output o_data_0_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[64] -----
	assign o_data_0_23_[0] = gfpga_pad_GPIO_PAD_fm[64];

// ----- Blif Benchmark output o_data_0_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[101] -----
	assign o_data_0_24_[0] = gfpga_pad_GPIO_PAD_fm[101];

// ----- Blif Benchmark output o_data_0_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[143] -----
	assign o_data_0_25_[0] = gfpga_pad_GPIO_PAD_fm[143];

// ----- Blif Benchmark output o_data_0_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[119] -----
	assign o_data_0_26_[0] = gfpga_pad_GPIO_PAD_fm[119];

// ----- Blif Benchmark output o_data_0_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[92] -----
	assign o_data_0_27_[0] = gfpga_pad_GPIO_PAD_fm[92];

// ----- Blif Benchmark output o_data_0_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[132] -----
	assign o_data_0_28_[0] = gfpga_pad_GPIO_PAD_fm[132];

// ----- Blif Benchmark output o_data_0_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[142] -----
	assign o_data_0_29_[0] = gfpga_pad_GPIO_PAD_fm[142];

// ----- Blif Benchmark output o_data_0_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[117] -----
	assign o_data_0_30_[0] = gfpga_pad_GPIO_PAD_fm[117];

// ----- Blif Benchmark output o_data_0_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[137] -----
	assign o_data_0_31_[0] = gfpga_pad_GPIO_PAD_fm[137];

// ----- Blif Benchmark output o_data_0_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[32] -----
	assign o_data_0_32_[0] = gfpga_pad_GPIO_PAD_fm[32];

// ----- Blif Benchmark output o_data_0_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[127] -----
	assign o_data_0_33_[0] = gfpga_pad_GPIO_PAD_fm[127];

// ----- Blif Benchmark output o_data_0_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[100] -----
	assign o_data_0_34_[0] = gfpga_pad_GPIO_PAD_fm[100];

// ----- Blif Benchmark output o_valid_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[34] -----
	assign o_valid_0[0] = gfpga_pad_GPIO_PAD_fm[34];

// ----- Blif Benchmark output o_vch_0 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[120] -----
	assign o_vch_0[0] = gfpga_pad_GPIO_PAD_fm[120];

// ----- Blif Benchmark output o_ack_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[108] -----
	assign o_ack_0_0_[0] = gfpga_pad_GPIO_PAD_fm[108];

// ----- Blif Benchmark output o_ack_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[83] -----
	assign o_ack_0_1_[0] = gfpga_pad_GPIO_PAD_fm[83];

// ----- Blif Benchmark output o_lck_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[110] -----
	assign o_lck_0_0_[0] = gfpga_pad_GPIO_PAD_fm[110];

// ----- Blif Benchmark output o_lck_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[90] -----
	assign o_lck_0_1_[0] = gfpga_pad_GPIO_PAD_fm[90];

// ----- Blif Benchmark output o_rdy_0_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[82] -----
	assign o_rdy_0_0_[0] = gfpga_pad_GPIO_PAD_fm[82];

// ----- Blif Benchmark output o_rdy_0_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[97] -----
	assign o_rdy_0_1_[0] = gfpga_pad_GPIO_PAD_fm[97];

// ----- Blif Benchmark output o_data_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[186] -----
	assign o_data_1_0_[0] = gfpga_pad_GPIO_PAD_fm[186];

// ----- Blif Benchmark output o_data_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[145] -----
	assign o_data_1_1_[0] = gfpga_pad_GPIO_PAD_fm[145];

// ----- Blif Benchmark output o_data_1_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[188] -----
	assign o_data_1_2_[0] = gfpga_pad_GPIO_PAD_fm[188];

// ----- Blif Benchmark output o_data_1_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[152] -----
	assign o_data_1_3_[0] = gfpga_pad_GPIO_PAD_fm[152];

// ----- Blif Benchmark output o_data_1_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[169] -----
	assign o_data_1_4_[0] = gfpga_pad_GPIO_PAD_fm[169];

// ----- Blif Benchmark output o_data_1_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[181] -----
	assign o_data_1_5_[0] = gfpga_pad_GPIO_PAD_fm[181];

// ----- Blif Benchmark output o_data_1_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[176] -----
	assign o_data_1_6_[0] = gfpga_pad_GPIO_PAD_fm[176];

// ----- Blif Benchmark output o_data_1_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[164] -----
	assign o_data_1_7_[0] = gfpga_pad_GPIO_PAD_fm[164];

// ----- Blif Benchmark output o_data_1_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[148] -----
	assign o_data_1_8_[0] = gfpga_pad_GPIO_PAD_fm[148];

// ----- Blif Benchmark output o_data_1_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[172] -----
	assign o_data_1_9_[0] = gfpga_pad_GPIO_PAD_fm[172];

// ----- Blif Benchmark output o_data_1_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[179] -----
	assign o_data_1_10_[0] = gfpga_pad_GPIO_PAD_fm[179];

// ----- Blif Benchmark output o_data_1_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[149] -----
	assign o_data_1_11_[0] = gfpga_pad_GPIO_PAD_fm[149];

// ----- Blif Benchmark output o_data_1_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[177] -----
	assign o_data_1_12_[0] = gfpga_pad_GPIO_PAD_fm[177];

// ----- Blif Benchmark output o_data_1_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[165] -----
	assign o_data_1_13_[0] = gfpga_pad_GPIO_PAD_fm[165];

// ----- Blif Benchmark output o_data_1_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[157] -----
	assign o_data_1_14_[0] = gfpga_pad_GPIO_PAD_fm[157];

// ----- Blif Benchmark output o_data_1_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[174] -----
	assign o_data_1_15_[0] = gfpga_pad_GPIO_PAD_fm[174];

// ----- Blif Benchmark output o_data_1_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[173] -----
	assign o_data_1_16_[0] = gfpga_pad_GPIO_PAD_fm[173];

// ----- Blif Benchmark output o_data_1_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[158] -----
	assign o_data_1_17_[0] = gfpga_pad_GPIO_PAD_fm[158];

// ----- Blif Benchmark output o_data_1_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[175] -----
	assign o_data_1_18_[0] = gfpga_pad_GPIO_PAD_fm[175];

// ----- Blif Benchmark output o_data_1_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[153] -----
	assign o_data_1_19_[0] = gfpga_pad_GPIO_PAD_fm[153];

// ----- Blif Benchmark output o_data_1_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[191] -----
	assign o_data_1_20_[0] = gfpga_pad_GPIO_PAD_fm[191];

// ----- Blif Benchmark output o_data_1_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[155] -----
	assign o_data_1_21_[0] = gfpga_pad_GPIO_PAD_fm[155];

// ----- Blif Benchmark output o_data_1_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[154] -----
	assign o_data_1_22_[0] = gfpga_pad_GPIO_PAD_fm[154];

// ----- Blif Benchmark output o_data_1_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[180] -----
	assign o_data_1_23_[0] = gfpga_pad_GPIO_PAD_fm[180];

// ----- Blif Benchmark output o_data_1_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[182] -----
	assign o_data_1_24_[0] = gfpga_pad_GPIO_PAD_fm[182];

// ----- Blif Benchmark output o_data_1_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[184] -----
	assign o_data_1_25_[0] = gfpga_pad_GPIO_PAD_fm[184];

// ----- Blif Benchmark output o_data_1_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[144] -----
	assign o_data_1_26_[0] = gfpga_pad_GPIO_PAD_fm[144];

// ----- Blif Benchmark output o_data_1_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[162] -----
	assign o_data_1_27_[0] = gfpga_pad_GPIO_PAD_fm[162];

// ----- Blif Benchmark output o_data_1_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[190] -----
	assign o_data_1_28_[0] = gfpga_pad_GPIO_PAD_fm[190];

// ----- Blif Benchmark output o_data_1_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[159] -----
	assign o_data_1_29_[0] = gfpga_pad_GPIO_PAD_fm[159];

// ----- Blif Benchmark output o_data_1_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[156] -----
	assign o_data_1_30_[0] = gfpga_pad_GPIO_PAD_fm[156];

// ----- Blif Benchmark output o_data_1_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[150] -----
	assign o_data_1_31_[0] = gfpga_pad_GPIO_PAD_fm[150];

// ----- Blif Benchmark output o_data_1_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[168] -----
	assign o_data_1_32_[0] = gfpga_pad_GPIO_PAD_fm[168];

// ----- Blif Benchmark output o_data_1_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[187] -----
	assign o_data_1_33_[0] = gfpga_pad_GPIO_PAD_fm[187];

// ----- Blif Benchmark output o_data_1_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[170] -----
	assign o_data_1_34_[0] = gfpga_pad_GPIO_PAD_fm[170];

// ----- Blif Benchmark output o_valid_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[178] -----
	assign o_valid_1[0] = gfpga_pad_GPIO_PAD_fm[178];

// ----- Blif Benchmark output o_vch_1 is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[166] -----
	assign o_vch_1[0] = gfpga_pad_GPIO_PAD_fm[166];

// ----- Blif Benchmark output o_ack_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[197] -----
	assign o_ack_1_0_[0] = gfpga_pad_GPIO_PAD_fm[197];

// ----- Blif Benchmark output o_ack_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[147] -----
	assign o_ack_1_1_[0] = gfpga_pad_GPIO_PAD_fm[147];

// ----- Blif Benchmark output o_lck_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[189] -----
	assign o_lck_1_0_[0] = gfpga_pad_GPIO_PAD_fm[189];

// ----- Blif Benchmark output o_lck_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[171] -----
	assign o_lck_1_1_[0] = gfpga_pad_GPIO_PAD_fm[171];

// ----- Blif Benchmark output o_rdy_1_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[183] -----
	assign o_rdy_1_0_[0] = gfpga_pad_GPIO_PAD_fm[183];

// ----- Blif Benchmark output o_rdy_1_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[185] -----
	assign o_rdy_1_1_[0] = gfpga_pad_GPIO_PAD_fm[185];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[33] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[35] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[40] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[41] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[42] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[44] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[47] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[48] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[50] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[53] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[54] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[55] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[63] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[69] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_5__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_6__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_7__8_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_8__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_7__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_6__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_5__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__0_.mem_top_track_34.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_34.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_0__0_.mem_top_track_52.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_0__0_.mem_top_track_52.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_out[0:7] = 8'b10000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_outb[0:7] = 8'b01111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_0__6_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__6_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__6_.mem_top_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__6_.mem_top_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__6_.mem_top_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__6_.mem_top_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__6_.mem_top_track_40.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__6_.mem_top_track_40.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__6_.mem_top_track_48.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__6_.mem_top_track_48.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__6_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__6_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__6_.mem_top_track_64.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_0__6_.mem_top_track_64.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_52.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_52.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__7_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_10.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_10.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_14.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_24.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_24.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_28.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_28.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_36.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_36.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_right_track_64.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_right_track_64.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_25.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_37.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_37.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_39.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_39.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_45.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_45.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_63.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_63.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_out[0:7] = 8'b00000010;
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_outb[0:7] = 8'b11111101;
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:9] = 10'b0001010000;
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:9] = 10'b1110101111;
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_out[0:9] = 10'b0001010000;
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_outb[0:9] = 10'b1110101111;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:9] = 10'b0001000010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:9] = 10'b1110111101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:9] = 10'b0001010000;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:9] = 10'b1110101111;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:9] = 10'b0001010000;
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:9] = 10'b1110101111;
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_right_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_1__7_.mem_right_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__7_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_15.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_15.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_49.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_49.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_left_track_17.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_1__7_.mem_left_track_17.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_1__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_left_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_left_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__7_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__7_.mem_left_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_left_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:5] = 6'b000010;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:5] = 6'b111101;
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_24.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__6_.mem_top_track_24.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__6_.mem_top_track_32.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_2__6_.mem_top_track_32.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_2__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_top_track_64.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_top_track_64.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_right_track_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__7_.mem_right_track_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_right_track_32.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_2__7_.mem_right_track_32.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_2__7_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__7_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_7.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_7.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_left_track_33.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_2__7_.mem_left_track_33.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_2__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__7_.mem_left_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_2__7_.mem_left_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_2__7_.mem_left_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_left_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_right_track_32.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_3__7_.mem_right_track_32.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_3__7_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_33.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_41.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_41.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_left_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_left_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_3__7_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_3__7_.mem_left_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_left_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_3__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_3__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__0_.mem_top_track_18.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_4__0_.mem_top_track_18.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_36.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_36.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_54.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_54.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_4__0_.mem_right_track_0.mem_out[0:9] = 10'b0000100100;
	force U0_formal_verification.sb_4__0_.mem_right_track_0.mem_outb[0:9] = 10'b1111011011;
	force U0_formal_verification.sb_4__0_.mem_right_track_8.mem_out[0:9] = 10'b0100000100;
	force U0_formal_verification.sb_4__0_.mem_right_track_8.mem_outb[0:9] = 10'b1011111011;
	force U0_formal_verification.sb_4__0_.mem_right_track_16.mem_out[0:7] = 8'b10000001;
	force U0_formal_verification.sb_4__0_.mem_right_track_16.mem_outb[0:7] = 8'b01111110;
	force U0_formal_verification.sb_4__0_.mem_right_track_24.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_4__0_.mem_right_track_24.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_4__0_.mem_right_track_32.mem_out[0:9] = 10'b0001000100;
	force U0_formal_verification.sb_4__0_.mem_right_track_32.mem_outb[0:9] = 10'b1110111011;
	force U0_formal_verification.sb_4__0_.mem_right_track_40.mem_out[0:9] = 10'b0001000100;
	force U0_formal_verification.sb_4__0_.mem_right_track_40.mem_outb[0:9] = 10'b1110111011;
	force U0_formal_verification.sb_4__0_.mem_right_track_48.mem_out[0:9] = 10'b0100000100;
	force U0_formal_verification.sb_4__0_.mem_right_track_48.mem_outb[0:9] = 10'b1011111011;
	force U0_formal_verification.sb_4__0_.mem_right_track_56.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_4__0_.mem_right_track_56.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_4__0_.mem_right_track_64.mem_out[0:9] = 10'b1000000100;
	force U0_formal_verification.sb_4__0_.mem_right_track_64.mem_outb[0:9] = 10'b0111111011;
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_4__1_.mem_right_track_0.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_4__1_.mem_right_track_0.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_4__1_.mem_right_track_8.mem_out[0:9] = 10'b0000100100;
	force U0_formal_verification.sb_4__1_.mem_right_track_8.mem_outb[0:9] = 10'b1111011011;
	force U0_formal_verification.sb_4__1_.mem_right_track_16.mem_out[0:9] = 10'b1000000100;
	force U0_formal_verification.sb_4__1_.mem_right_track_16.mem_outb[0:9] = 10'b0111111011;
	force U0_formal_verification.sb_4__1_.mem_right_track_24.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_4__1_.mem_right_track_24.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_4__1_.mem_right_track_32.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_4__1_.mem_right_track_32.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_4__1_.mem_right_track_40.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_4__1_.mem_right_track_40.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_4__1_.mem_right_track_48.mem_out[0:7] = 8'b10000001;
	force U0_formal_verification.sb_4__1_.mem_right_track_48.mem_outb[0:7] = 8'b01111110;
	force U0_formal_verification.sb_4__1_.mem_right_track_56.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_4__1_.mem_right_track_56.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_4__1_.mem_right_track_64.mem_out[0:9] = 10'b0100000100;
	force U0_formal_verification.sb_4__1_.mem_right_track_64.mem_outb[0:9] = 10'b1011111011;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:9] = 10'b1000000010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_outb[0:9] = 10'b0111111101;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_out[0:9] = 10'b0000100100;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_outb[0:9] = 10'b1111011011;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_out[0:9] = 10'b0100000010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_outb[0:9] = 10'b1011111101;
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__2_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__2_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__2_.mem_right_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__2_.mem_right_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__2_.mem_right_track_16.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_4__2_.mem_right_track_16.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_4__2_.mem_right_track_24.mem_out[0:7] = 8'b00000010;
	force U0_formal_verification.sb_4__2_.mem_right_track_24.mem_outb[0:7] = 8'b11111101;
	force U0_formal_verification.sb_4__2_.mem_right_track_32.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_4__2_.mem_right_track_32.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_4__2_.mem_right_track_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_4__2_.mem_right_track_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_4__2_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__2_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__2_.mem_right_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__2_.mem_right_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__2_.mem_right_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__2_.mem_right_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:7] = 8'b00000010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_right_track_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__3_.mem_right_track_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__3_.mem_right_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__3_.mem_right_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__3_.mem_right_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__3_.mem_right_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__3_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__3_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__3_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_right_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__3_.mem_right_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__3_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__3_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__3_.mem_right_track_56.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__3_.mem_right_track_56.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__3_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__3_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__4_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__4_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__4_.mem_right_track_8.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__4_.mem_right_track_8.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__4_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_right_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__4_.mem_right_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__4_.mem_right_track_32.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__4_.mem_right_track_32.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__4_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_right_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__4_.mem_right_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__4_.mem_right_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__4_.mem_right_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__4_.mem_right_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__4_.mem_right_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__5_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_right_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__5_.mem_right_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__5_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__5_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__6_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_right_track_24.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__6_.mem_right_track_24.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_4__7_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_4__7_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_23.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_23.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_33.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_left_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_left_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_4__7_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_4__7_.mem_left_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_left_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_4__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_4__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_4.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_5__0_.mem_top_track_4.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_5__0_.mem_top_track_6.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__0_.mem_top_track_6.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__0_.mem_top_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__0_.mem_top_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__0_.mem_top_track_10.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_top_track_10.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_top_track_12.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_12.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_14.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__0_.mem_top_track_14.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__0_.mem_top_track_16.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__0_.mem_top_track_16.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__0_.mem_top_track_18.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_18.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_20.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_5__0_.mem_top_track_20.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_5__0_.mem_top_track_22.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_5__0_.mem_top_track_22.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_5__0_.mem_top_track_24.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__0_.mem_top_track_24.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__0_.mem_top_track_26.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__0_.mem_top_track_26.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__0_.mem_top_track_28.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__0_.mem_top_track_28.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__0_.mem_top_track_30.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_top_track_30.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_top_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_34.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_5__0_.mem_top_track_34.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_5__0_.mem_top_track_36.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_36.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_38.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_5__0_.mem_top_track_38.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_5__0_.mem_top_track_40.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_top_track_40.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_top_track_42.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_42.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_44.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_44.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_46.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_46.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_top_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_top_track_50.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_5__0_.mem_top_track_50.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_5__0_.mem_top_track_52.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.sb_5__0_.mem_top_track_52.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.sb_5__0_.mem_top_track_54.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_54.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_top_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__0_.mem_top_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__0_.mem_top_track_58.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_top_track_58.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_top_track_60.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__0_.mem_top_track_60.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__0_.mem_top_track_62.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__0_.mem_top_track_62.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__0_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__0_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__0_.mem_right_track_0.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__0_.mem_right_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__0_.mem_right_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__0_.mem_right_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__0_.mem_right_track_16.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__0_.mem_right_track_16.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__0_.mem_right_track_24.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__0_.mem_right_track_24.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__0_.mem_right_track_32.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__0_.mem_right_track_32.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__0_.mem_right_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__0_.mem_right_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__0_.mem_right_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__0_.mem_right_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__0_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__0_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__0_.mem_right_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__0_.mem_right_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__0_.mem_left_track_1.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__0_.mem_left_track_1.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__0_.mem_left_track_9.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_5__0_.mem_left_track_9.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_5__0_.mem_left_track_17.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_5__0_.mem_left_track_17.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_5__0_.mem_left_track_25.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_5__0_.mem_left_track_25.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_5__0_.mem_left_track_33.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_5__0_.mem_left_track_33.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_5__0_.mem_left_track_41.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__0_.mem_left_track_41.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__0_.mem_left_track_49.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_5__0_.mem_left_track_49.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_5__0_.mem_left_track_57.mem_out[0:7] = 8'b10000001;
	force U0_formal_verification.sb_5__0_.mem_left_track_57.mem_outb[0:7] = 8'b01111110;
	force U0_formal_verification.sb_5__0_.mem_left_track_65.mem_out[0:9] = 10'b0100000010;
	force U0_formal_verification.sb_5__0_.mem_left_track_65.mem_outb[0:9] = 10'b1011111101;
	force U0_formal_verification.sb_5__1_.mem_top_track_0.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_5__1_.mem_top_track_0.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_5__1_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__1_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__1_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__1_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__1_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__1_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__1_.mem_top_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__1_.mem_top_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__1_.mem_top_track_40.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_5__1_.mem_top_track_40.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_5__1_.mem_top_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__1_.mem_top_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__1_.mem_top_track_56.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__1_.mem_top_track_56.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__1_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__1_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__1_.mem_right_track_0.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__1_.mem_right_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__1_.mem_right_track_8.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__1_.mem_right_track_8.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__1_.mem_right_track_16.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_5__1_.mem_right_track_16.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_5__1_.mem_right_track_24.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_5__1_.mem_right_track_24.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_5__1_.mem_right_track_32.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_5__1_.mem_right_track_32.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_5__1_.mem_right_track_40.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__1_.mem_right_track_40.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__1_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__1_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__1_.mem_right_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__1_.mem_right_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__1_.mem_right_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__1_.mem_right_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_out[0:9] = 10'b1000010000;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_17.mem_outb[0:9] = 10'b0111101111;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_out[0:9] = 10'b0001000010;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_25.mem_outb[0:9] = 10'b1110111101;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_out[0:9] = 10'b0010000100;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_33.mem_outb[0:9] = 10'b1101111011;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_41.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_41.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_49.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_49.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_57.mem_out[0:9] = 10'b0001010000;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_57.mem_outb[0:9] = 10'b1110101111;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_65.mem_out[0:9] = 10'b0001000010;
	force U0_formal_verification.sb_5__1_.mem_bottom_track_65.mem_outb[0:9] = 10'b1110111101;
	force U0_formal_verification.sb_5__1_.mem_left_track_1.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__1_.mem_left_track_1.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__1_.mem_left_track_9.mem_out[0:9] = 10'b0010010000;
	force U0_formal_verification.sb_5__1_.mem_left_track_9.mem_outb[0:9] = 10'b1101101111;
	force U0_formal_verification.sb_5__1_.mem_left_track_17.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_5__1_.mem_left_track_17.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_5__1_.mem_left_track_25.mem_out[0:9] = 10'b0100001000;
	force U0_formal_verification.sb_5__1_.mem_left_track_25.mem_outb[0:9] = 10'b1011110111;
	force U0_formal_verification.sb_5__1_.mem_left_track_33.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__1_.mem_left_track_33.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__1_.mem_left_track_41.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__1_.mem_left_track_41.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__1_.mem_left_track_49.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_5__1_.mem_left_track_49.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_5__1_.mem_left_track_57.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.sb_5__1_.mem_left_track_57.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.sb_5__1_.mem_left_track_65.mem_out[0:9] = 10'b0010000010;
	force U0_formal_verification.sb_5__1_.mem_left_track_65.mem_outb[0:9] = 10'b1101111101;
	force U0_formal_verification.sb_5__2_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__2_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__2_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__2_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__2_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__2_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__2_.mem_top_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__2_.mem_top_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__2_.mem_top_track_32.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__2_.mem_top_track_32.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__2_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__2_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__2_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__2_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__2_.mem_top_track_56.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__2_.mem_top_track_56.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__2_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__2_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__2_.mem_right_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__2_.mem_right_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__2_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__2_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__2_.mem_right_track_16.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_5__2_.mem_right_track_16.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_5__2_.mem_right_track_24.mem_out[0:7] = 8'b00000010;
	force U0_formal_verification.sb_5__2_.mem_right_track_24.mem_outb[0:7] = 8'b11111101;
	force U0_formal_verification.sb_5__2_.mem_right_track_32.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_5__2_.mem_right_track_32.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_5__2_.mem_right_track_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_5__2_.mem_right_track_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_5__2_.mem_right_track_48.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__2_.mem_right_track_48.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__2_.mem_right_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__2_.mem_right_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__2_.mem_right_track_64.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__2_.mem_right_track_64.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_out[0:7] = 8'b00000010;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b11111101;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_41.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_57.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_65.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_5__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_5__2_.mem_left_track_1.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.sb_5__2_.mem_left_track_1.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_5__2_.mem_left_track_9.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__2_.mem_left_track_9.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__2_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__2_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__2_.mem_left_track_25.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__2_.mem_left_track_25.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__2_.mem_left_track_33.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_5__2_.mem_left_track_33.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_5__2_.mem_left_track_41.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.sb_5__2_.mem_left_track_41.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.sb_5__2_.mem_left_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__2_.mem_left_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__2_.mem_left_track_57.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__2_.mem_left_track_57.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__2_.mem_left_track_65.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__2_.mem_left_track_65.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_top_track_24.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_top_track_24.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__3_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__3_.mem_right_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__3_.mem_right_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__3_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_right_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__3_.mem_right_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__3_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_right_track_40.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__3_.mem_right_track_40.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__3_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_right_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__3_.mem_right_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_41.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_49.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_left_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__3_.mem_left_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__3_.mem_left_track_9.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__3_.mem_left_track_9.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__3_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_left_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_left_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_left_track_33.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__3_.mem_left_track_33.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__3_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__3_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__3_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__3_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__3_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__3_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__3_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__3_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__4_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__4_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__4_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__4_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__4_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__4_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__4_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_top_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_top_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_top_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__4_.mem_top_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__4_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__4_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__4_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_right_track_16.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__4_.mem_right_track_16.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__4_.mem_right_track_24.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_right_track_24.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__4_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__4_.mem_right_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_right_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__4_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__4_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_right_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__4_.mem_right_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_65.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_left_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_5__4_.mem_left_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_5__4_.mem_left_track_9.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_left_track_9.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__4_.mem_left_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_5__4_.mem_left_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_5__4_.mem_left_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__4_.mem_left_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__4_.mem_left_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__4_.mem_left_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__4_.mem_left_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__4_.mem_left_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__4_.mem_left_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__4_.mem_left_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__4_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__4_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__5_.mem_top_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__5_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_right_track_40.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__5_.mem_right_track_40.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__5_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__5_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__5_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__5_.mem_left_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__5_.mem_left_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__5_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__5_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__5_.mem_left_track_49.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__5_.mem_left_track_49.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__5_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__5_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__5_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__6_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_5__6_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_5__6_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_5__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_5__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__7_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_5__7_.mem_left_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_left_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_5__7_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_5__7_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_5__7_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_5__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_5__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__0_.mem_top_track_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__0_.mem_top_track_2.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_32.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_34.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__0_.mem_top_track_34.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__0_.mem_top_track_36.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__0_.mem_top_track_36.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__0_.mem_top_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_6__0_.mem_top_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_6__0_.mem_top_track_52.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_62.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_64.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__0_.mem_top_track_64.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__0_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__0_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__0_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__0_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__0_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__0_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__0_.mem_right_track_24.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__0_.mem_right_track_24.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__0_.mem_right_track_32.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__0_.mem_right_track_32.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__0_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__0_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__0_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__0_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__0_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__0_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__0_.mem_right_track_64.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__0_.mem_right_track_64.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__0_.mem_left_track_1.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__0_.mem_left_track_1.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__0_.mem_left_track_9.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__0_.mem_left_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__0_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__0_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__0_.mem_left_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__0_.mem_left_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__0_.mem_left_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__0_.mem_left_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__0_.mem_left_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__0_.mem_left_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__0_.mem_left_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__0_.mem_left_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__0_.mem_left_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__0_.mem_left_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__0_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__0_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__1_.mem_top_track_0.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_6__1_.mem_top_track_0.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_6__1_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__1_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__1_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__1_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__1_.mem_top_track_24.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__1_.mem_top_track_24.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__1_.mem_top_track_32.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.sb_6__1_.mem_top_track_32.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.sb_6__1_.mem_top_track_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_6__1_.mem_top_track_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_6__1_.mem_top_track_48.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__1_.mem_top_track_48.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__1_.mem_top_track_56.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__1_.mem_top_track_56.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__1_.mem_top_track_64.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__1_.mem_top_track_64.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__1_.mem_right_track_0.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__1_.mem_right_track_0.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__1_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__1_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__1_.mem_right_track_16.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.sb_6__1_.mem_right_track_16.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.sb_6__1_.mem_right_track_24.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__1_.mem_right_track_24.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__1_.mem_right_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__1_.mem_right_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__1_.mem_right_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__1_.mem_right_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__1_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__1_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__1_.mem_right_track_56.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__1_.mem_right_track_56.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__1_.mem_right_track_64.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__1_.mem_right_track_64.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__1_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__1_.mem_left_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__1_.mem_left_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__1_.mem_left_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__1_.mem_left_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__1_.mem_left_track_17.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__1_.mem_left_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__1_.mem_left_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__1_.mem_left_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__1_.mem_left_track_33.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_6__1_.mem_left_track_33.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_6__1_.mem_left_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__1_.mem_left_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__1_.mem_left_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__1_.mem_left_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__1_.mem_left_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__1_.mem_left_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__1_.mem_left_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__1_.mem_left_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__2_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__2_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__2_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__2_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__2_.mem_top_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__2_.mem_top_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__2_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__2_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__2_.mem_top_track_48.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__2_.mem_top_track_48.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__2_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__2_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__2_.mem_top_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__2_.mem_top_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__2_.mem_right_track_0.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__2_.mem_right_track_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__2_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_right_track_16.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_6__2_.mem_right_track_16.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_6__2_.mem_right_track_24.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__2_.mem_right_track_24.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__2_.mem_right_track_32.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__2_.mem_right_track_32.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__2_.mem_right_track_40.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_6__2_.mem_right_track_40.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_6__2_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__2_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__2_.mem_right_track_64.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__2_.mem_right_track_64.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_17.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_25.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_33.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_41.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_41.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_57.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_65.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_6__2_.mem_bottom_track_65.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_6__2_.mem_left_track_1.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_6__2_.mem_left_track_1.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_6__2_.mem_left_track_9.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__2_.mem_left_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__2_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__2_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__2_.mem_left_track_25.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__2_.mem_left_track_25.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__2_.mem_left_track_33.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.sb_6__2_.mem_left_track_33.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.sb_6__2_.mem_left_track_41.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.sb_6__2_.mem_left_track_41.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_6__2_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__2_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__2_.mem_left_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__2_.mem_left_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__2_.mem_left_track_65.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__2_.mem_left_track_65.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__3_.mem_top_track_0.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__3_.mem_top_track_0.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__3_.mem_top_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__3_.mem_top_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__3_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_top_track_48.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__3_.mem_top_track_48.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__3_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_top_track_64.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_top_track_64.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_right_track_0.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_right_track_0.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_right_track_8.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__3_.mem_right_track_8.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__3_.mem_right_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__3_.mem_right_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__3_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__3_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_41.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_57.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__3_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__3_.mem_left_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_left_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_left_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__3_.mem_left_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__3_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__3_.mem_left_track_33.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__3_.mem_left_track_33.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__3_.mem_left_track_41.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__3_.mem_left_track_41.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__3_.mem_left_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__3_.mem_left_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__3_.mem_left_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__3_.mem_left_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__3_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__3_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__4_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__4_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_right_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__4_.mem_right_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__4_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_right_track_48.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__4_.mem_right_track_48.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__4_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_right_track_64.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__4_.mem_right_track_64.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_57.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_left_track_9.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__4_.mem_left_track_9.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__4_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_left_track_25.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__4_.mem_left_track_25.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__4_.mem_left_track_33.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__4_.mem_left_track_33.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__4_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__4_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__4_.mem_left_track_49.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__4_.mem_left_track_49.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__4_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__4_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__4_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_top_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__5_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__5_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_right_track_48.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__5_.mem_right_track_48.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__5_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__5_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_41.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_49.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_left_track_25.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__5_.mem_left_track_25.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__5_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__5_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__5_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__5_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__5_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_24.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_top_track_24.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_top_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_top_track_56.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__6_.mem_top_track_56.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__6_.mem_top_track_64.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_top_track_64.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__6_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__6_.mem_right_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_right_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_24.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_right_track_24.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_32.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_right_track_32.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_40.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_right_track_40.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_48.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_right_track_48.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_right_track_56.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_right_track_56.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__6_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_1.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_1.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_25.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_25.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_33.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_left_track_33.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_left_track_41.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_left_track_41.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_left_track_49.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_6__6_.mem_left_track_49.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_6__6_.mem_left_track_57.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_57.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__6_.mem_left_track_65.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__6_.mem_left_track_65.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_right_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_right_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_right_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_right_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_right_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_right_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_right_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_right_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_right_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_right_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_right_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_right_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_right_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_right_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_6__7_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_left_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_left_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_left_track_17.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_6__7_.mem_left_track_17.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_6__7_.mem_left_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_left_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_left_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_left_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_left_track_41.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_left_track_41.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_left_track_49.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_6__7_.mem_left_track_49.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_6__7_.mem_left_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_left_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_6__7_.mem_left_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_6__7_.mem_left_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__0_.mem_top_track_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_2.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_2.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_6.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_8.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_8.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_14.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_14.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_18.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_18.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_32.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_32.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_34.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_34.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_38.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_38.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_42.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_42.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_48.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_48.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_50.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_56.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_56.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_58.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_top_track_58.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_1.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_3.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_9.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_11.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_15.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_19.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_19.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_23.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_left_track_23.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_left_track_25.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_25.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_27.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_27.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_33.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_33.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_35.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_35.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_37.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_37.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_45.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__0_.mem_left_track_45.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__0_.mem_left_track_47.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_47.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_49.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_49.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_51.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_51.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_57.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_57.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_59.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_59.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_top_track_0.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_7__1_.mem_top_track_0.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_7__1_.mem_top_track_8.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__1_.mem_top_track_8.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__1_.mem_top_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__1_.mem_top_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__1_.mem_top_track_24.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__1_.mem_top_track_24.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__1_.mem_top_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__1_.mem_top_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__1_.mem_top_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__1_.mem_top_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__1_.mem_top_track_48.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__1_.mem_top_track_48.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__1_.mem_top_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__1_.mem_top_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__1_.mem_top_track_64.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__1_.mem_top_track_64.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_33.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_49.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_49.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_65.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__1_.mem_bottom_track_65.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__1_.mem_left_track_1.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_3.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_3.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_5.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_5.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_11.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_11.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_33.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_33.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_35.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_35.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_49.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__1_.mem_left_track_49.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__1_.mem_left_track_51.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_51.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_59.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__1_.mem_left_track_59.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__1_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__1_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_top_track_0.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__2_.mem_top_track_0.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__2_.mem_top_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__2_.mem_top_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__2_.mem_top_track_16.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__2_.mem_top_track_16.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__2_.mem_top_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__2_.mem_top_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__2_.mem_top_track_32.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__2_.mem_top_track_32.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__2_.mem_top_track_40.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__2_.mem_top_track_40.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__2_.mem_top_track_48.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__2_.mem_top_track_48.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__2_.mem_top_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__2_.mem_top_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__2_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__2_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_9.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_25.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_49.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_49.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_57.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_57.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_65.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__2_.mem_bottom_track_65.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__2_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__2_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__2_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_7.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__2_.mem_left_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__2_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_25.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_25.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__2_.mem_left_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__2_.mem_left_track_29.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_29.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_39.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__2_.mem_left_track_39.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__2_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_43.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_43.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_47.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__2_.mem_left_track_47.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__2_.mem_left_track_49.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__2_.mem_left_track_49.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__2_.mem_left_track_51.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__2_.mem_left_track_51.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__2_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_57.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__2_.mem_left_track_57.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__2_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__2_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__3_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__3_.mem_top_track_8.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__3_.mem_top_track_8.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__3_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__3_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__3_.mem_top_track_24.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__3_.mem_top_track_24.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__3_.mem_top_track_32.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__3_.mem_top_track_32.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__3_.mem_top_track_40.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__3_.mem_top_track_40.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__3_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__3_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__3_.mem_top_track_56.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__3_.mem_top_track_56.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__3_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__3_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_17.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_25.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_33.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_41.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_41.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_49.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_49.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_57.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_57.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_65.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_65.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__3_.mem_left_track_1.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__3_.mem_left_track_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__3_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_7.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_9.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_15.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__3_.mem_left_track_15.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__3_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_23.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_23.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__3_.mem_left_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_33.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__3_.mem_left_track_33.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__3_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_51.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_51.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__3_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__4_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__4_.mem_top_track_8.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__4_.mem_top_track_8.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__4_.mem_top_track_16.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__4_.mem_top_track_16.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__4_.mem_top_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__4_.mem_top_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__4_.mem_top_track_32.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__4_.mem_top_track_32.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__4_.mem_top_track_40.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__4_.mem_top_track_40.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__4_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__4_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__4_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__4_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__4_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__4_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_9.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_17.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_25.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_out[0:5] = 6'b100001;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_33.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_41.mem_out[0:5] = 6'b100010;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_41.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_49.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_49.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__4_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__4_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_11.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__4_.mem_left_track_11.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__4_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_21.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__4_.mem_left_track_21.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__4_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_41.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__4_.mem_left_track_41.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__4_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_61.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_61.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__4_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__5_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__5_.mem_top_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_top_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_top_track_16.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_top_track_16.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_top_track_24.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__5_.mem_top_track_24.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__5_.mem_top_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__5_.mem_top_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__5_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__5_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__5_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__5_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__5_.mem_top_track_56.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__5_.mem_top_track_56.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__5_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_9.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_out[0:5] = 6'b001010;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_25.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_33.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_41.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_41.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_49.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_49.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_57.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_57.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__5_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_13.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__5_.mem_left_track_13.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__5_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_27.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__5_.mem_left_track_27.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__5_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_31.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_31.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_35.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__5_.mem_left_track_35.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__5_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_43.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__5_.mem_left_track_43.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__5_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_61.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__5_.mem_left_track_61.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__5_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__5_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_top_track_0.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_top_track_0.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_top_track_8.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_top_track_8.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_top_track_16.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_top_track_16.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_top_track_24.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_top_track_24.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_top_track_32.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_top_track_32.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_top_track_40.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_top_track_40.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_top_track_48.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_top_track_48.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_top_track_56.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_top_track_56.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_top_track_64.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_top_track_64.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_out[0:5] = 6'b010010;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_outb[0:5] = 6'b101101;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_9.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_17.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_25.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_33.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_41.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_41.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_49.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_49.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_57.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_57.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_65.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_7__6_.mem_bottom_track_65.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_7__6_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_35.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__6_.mem_left_track_35.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__6_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_49.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_7__6_.mem_left_track_49.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_7__6_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__6_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_29.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_41.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_41.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__7_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_16.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_16.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_17.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_17.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_18.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_18.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_19.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_19.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_20.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_20.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_21.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_21.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_22.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_22.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_23.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_23.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_24.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_24.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_25.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_25.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_26.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_26.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_27.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_27.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_28.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_28.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_29.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_29.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_30.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_30.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_31.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_31.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_32.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_32.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_33.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_33.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_34.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_34.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_35.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_35.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_36.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_36.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_37.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_37.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_38.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_38.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_39.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_39.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_40.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_40.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_41.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_41.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_42.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_42.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_43.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_43.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_44.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_44.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_45.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_45.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_46.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_46.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_47.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_47.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_48.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_48.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_49.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_49.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_50.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_50.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_51.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_51.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_8.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_8.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_9.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_9.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_10.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_10.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_11.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_11.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_12.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_12.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_13.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_13.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_14.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_14.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_15.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_15.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_16.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_16.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_17.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_17.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_18.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_18.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_19.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_19.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_20.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_20.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_21.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_21.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_22.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_22.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_23.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_23.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_24.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_24.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_25.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_25.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_26.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_26.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_27.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_27.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_28.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_28.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_29.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_29.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_30.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_30.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_31.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_31.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_32.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_32.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_33.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_33.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_34.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_34.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_35.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_35.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_36.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_36.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_37.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_37.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_38.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_38.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_39.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_39.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_40.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_40.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_41.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_41.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_42.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_42.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_43.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_43.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_44.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_44.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_45.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_45.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_46.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_46.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_47.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_47.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_48.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_48.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_49.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_49.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_50.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_50.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_51.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_51.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_52.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_52.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_1__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_2__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_3__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_4__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_1.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_2.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_4.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_5.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_6.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_8.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_9.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_10.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_10.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_11.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_11.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_12.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_12.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_13.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_13.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_14.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_14.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_15.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_15.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_16.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_16.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_17.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_17.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_18.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_18.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_19.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_19.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_20.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_20.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_21.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_21.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_22.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_22.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_23.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_23.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_24.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_24.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_25.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_25.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_26.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_26.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_27.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_27.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_28.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_28.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_29.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_29.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_30.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_30.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_31.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_31.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_32.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_32.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_33.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_33.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_34.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_34.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_35.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_35.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_36.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_36.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_37.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_37.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_38.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_38.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_39.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_39.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_40.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_40.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_41.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_41.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_42.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_42.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_43.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_43.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_44.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_44.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_45.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_45.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_46.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_46.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_47.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_47.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_48.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_48.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_49.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_49.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_50.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_50.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_51.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__0_.mem_bottom_ipin_51.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_8.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_8.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_9.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_9.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_10.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_10.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_11.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_11.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_12.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_12.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_13.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_13.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_14.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_14.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_15.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_15.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_16.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_16.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_17.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_17.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_18.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_18.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_19.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_19.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_20.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_20.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_21.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_21.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_22.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_22.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_23.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_23.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_24.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_24.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_25.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_25.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_26.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_26.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_27.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_27.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_28.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_28.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_29.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_29.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_30.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_30.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_31.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_31.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_32.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_32.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_33.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_33.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_34.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_34.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_35.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_35.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_36.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_36.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_37.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_37.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_38.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_38.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_39.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_39.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_40.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_40.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_41.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_41.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_42.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_42.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_43.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_43.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_44.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_44.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_45.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_45.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_46.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_46.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_47.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_47.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_48.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_48.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_49.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_49.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_50.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_50.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_51.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_51.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_52.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_52.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_5__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_6__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_5.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_7.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__1_.mem_bottom_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cbx_7__7_.mem_bottom_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_2.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_2.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_3.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_3.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_4.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_4.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_5.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_5.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_6.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_6.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_7.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_7.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_8.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_8.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_9.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_9.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_10.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_10.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_11.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_11.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_12.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_12.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_13.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_13.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_14.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_14.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_15.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_15.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_16.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_16.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_17.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_17.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_18.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_18.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_19.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_19.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_20.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_20.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_21.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_21.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_22.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_22.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_23.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_23.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_24.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_24.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_25.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_25.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_26.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_26.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_27.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_27.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_28.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_28.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_29.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_29.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_30.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_30.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_31.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_31.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_32.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_32.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_33.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_33.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_34.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_34.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_35.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_35.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_36.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_36.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_37.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_37.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_38.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_38.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_39.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_39.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_40.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_40.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_41.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_41.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_42.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_42.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_43.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_43.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_44.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_44.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_45.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_45.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_46.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_46.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_47.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_47.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_48.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_48.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_49.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_49.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_50.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_50.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_51.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_51.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_0__7_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_16.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_16.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_17.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_17.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_18.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_18.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_19.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_19.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_20.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_20.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_21.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_21.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_22.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_22.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_23.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_23.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_24.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_24.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_25.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_25.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_26.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_26.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_27.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_27.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_28.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_28.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_29.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_29.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_30.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_30.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_31.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_31.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_32.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_32.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_33.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_33.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_34.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_34.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_35.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_35.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_36.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_36.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_37.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_37.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_38.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_38.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_39.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_39.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_40.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_40.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_41.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_41.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_42.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_42.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_43.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_43.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_44.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_44.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_45.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_45.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_46.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_46.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_47.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_47.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_48.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_48.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_49.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_49.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_50.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_50.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_51.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_51.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_52.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_52.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_8.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_8.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_9.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_9.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_10.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_10.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_11.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_11.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_12.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_12.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_13.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_13.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_14.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_14.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_15.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_15.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_16.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_16.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_17.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_17.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_18.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_18.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_19.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_19.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_20.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_20.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_21.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_21.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_22.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_22.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_23.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_23.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_24.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_24.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_25.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_25.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_26.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_26.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_27.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_27.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_28.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_28.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_29.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_29.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_30.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_30.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_31.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_31.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_32.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_32.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_33.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_33.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_34.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_34.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_35.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_35.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_36.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_36.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_37.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_37.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_38.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_38.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_39.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_39.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_40.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_40.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_41.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_41.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_42.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_42.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_43.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_43.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_44.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_44.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_45.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_45.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_46.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_46.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_47.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_47.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_48.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_48.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_49.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_49.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_50.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_50.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_51.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_51.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_8.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_8.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_9.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_9.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_10.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_10.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_11.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_11.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_12.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_12.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_13.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_13.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_14.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_14.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_15.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_15.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_16.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_16.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_17.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_17.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_18.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_18.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_19.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_19.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_20.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_20.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_21.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_21.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_22.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_22.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_23.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_23.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_24.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_24.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_25.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_25.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_26.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_26.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_27.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_27.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_28.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_28.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_29.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_29.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_30.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_30.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_31.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_31.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_32.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_32.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_33.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_33.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_34.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_34.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_35.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_35.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_36.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_36.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_37.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_37.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_38.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_38.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_39.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_39.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_40.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_40.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_41.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_41.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_42.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_42.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_43.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_43.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_44.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_44.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_45.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_45.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_46.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_46.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_47.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_47.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_48.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_48.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_49.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_49.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_50.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_50.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_51.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_51.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_52.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_5__1_.mem_right_ipin_52.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_5__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_left_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_6__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_4.mem_out[0:7] = 8'b01000010;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_4.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_5.mem_out[0:7] = 8'b00100100;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_5.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_6.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_6.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_7.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_7__1_.mem_left_ipin_7.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_0.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_0.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_1.mem_out[0:7] = 8'b10000010;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_1.mem_outb[0:7] = 8'b01111101;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_3.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_3.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_4.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_4.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_5.mem_out[0:7] = 8'b00101000;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_5.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__2_.mem_right_ipin_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_0.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_0.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_1.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_1.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_2.mem_out[0:7] = 8'b00010010;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_2.mem_outb[0:7] = 8'b11101101;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_3.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_3.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_4.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_4.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_6.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_6.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__3_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_1.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_1.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_2.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_2.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_3.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_3.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_4.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_4.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_5.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_5.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_7.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_7__4_.mem_left_ipin_7.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_7.mem_out[0:7] = 8'b10001000;
	force U0_formal_verification.cby_7__5_.mem_left_ipin_7.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_0.mem_out[0:7] = 8'b01001000;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_0.mem_outb[0:7] = 8'b10110111;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_3.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_3.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_4.mem_out[0:7] = 8'b00100010;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_4.mem_outb[0:7] = 8'b11011101;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_6.mem_out[0:7] = 8'b10000100;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_6.mem_outb[0:7] = 8'b01111011;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__6_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_2.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_2.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_3.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_3.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_4.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_4.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_5.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_5.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_6.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_6.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_7.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.cby_7__7_.mem_left_ipin_7.mem_outb[0:7] = 8'b11111110;
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for mesh_bench_top_formal_verification -----

//----- Default net type -----
`default_nettype wire

