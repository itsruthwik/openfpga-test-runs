//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Sep 25 16:03:58 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(pReset,
                prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:703] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:228] cbx_1__0__0_chanx_left_out;
wire [0:228] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__10_ccff_tail;
wire [0:228] cbx_1__0__10_chanx_left_out;
wire [0:228] cbx_1__0__10_chanx_right_out;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__11_ccff_tail;
wire [0:228] cbx_1__0__11_chanx_left_out;
wire [0:228] cbx_1__0__11_chanx_right_out;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__12_ccff_tail;
wire [0:228] cbx_1__0__12_chanx_left_out;
wire [0:228] cbx_1__0__12_chanx_right_out;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__13_ccff_tail;
wire [0:228] cbx_1__0__13_chanx_left_out;
wire [0:228] cbx_1__0__13_chanx_right_out;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__14_ccff_tail;
wire [0:228] cbx_1__0__14_chanx_left_out;
wire [0:228] cbx_1__0__14_chanx_right_out;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__15_ccff_tail;
wire [0:228] cbx_1__0__15_chanx_left_out;
wire [0:228] cbx_1__0__15_chanx_right_out;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__16_ccff_tail;
wire [0:228] cbx_1__0__16_chanx_left_out;
wire [0:228] cbx_1__0__16_chanx_right_out;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__17_ccff_tail;
wire [0:228] cbx_1__0__17_chanx_left_out;
wire [0:228] cbx_1__0__17_chanx_right_out;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__18_ccff_tail;
wire [0:228] cbx_1__0__18_chanx_left_out;
wire [0:228] cbx_1__0__18_chanx_right_out;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__19_ccff_tail;
wire [0:228] cbx_1__0__19_chanx_left_out;
wire [0:228] cbx_1__0__19_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:228] cbx_1__0__1_chanx_left_out;
wire [0:228] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__20_ccff_tail;
wire [0:228] cbx_1__0__20_chanx_left_out;
wire [0:228] cbx_1__0__20_chanx_right_out;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__21_ccff_tail;
wire [0:228] cbx_1__0__21_chanx_left_out;
wire [0:228] cbx_1__0__21_chanx_right_out;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:228] cbx_1__0__2_chanx_left_out;
wire [0:228] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:228] cbx_1__0__3_chanx_left_out;
wire [0:228] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:228] cbx_1__0__4_chanx_left_out;
wire [0:228] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:228] cbx_1__0__5_chanx_left_out;
wire [0:228] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__6_ccff_tail;
wire [0:228] cbx_1__0__6_chanx_left_out;
wire [0:228] cbx_1__0__6_chanx_right_out;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__7_ccff_tail;
wire [0:228] cbx_1__0__7_chanx_left_out;
wire [0:228] cbx_1__0__7_chanx_right_out;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__8_ccff_tail;
wire [0:228] cbx_1__0__8_chanx_left_out;
wire [0:228] cbx_1__0__8_chanx_right_out;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__9_ccff_tail;
wire [0:228] cbx_1__0__9_chanx_left_out;
wire [0:228] cbx_1__0__9_chanx_right_out;
wire [0:228] cbx_1__1__0_chanx_left_out;
wire [0:228] cbx_1__1__0_chanx_right_out;
wire [0:228] cbx_1__1__100_chanx_left_out;
wire [0:228] cbx_1__1__100_chanx_right_out;
wire [0:228] cbx_1__1__101_chanx_left_out;
wire [0:228] cbx_1__1__101_chanx_right_out;
wire [0:228] cbx_1__1__102_chanx_left_out;
wire [0:228] cbx_1__1__102_chanx_right_out;
wire [0:228] cbx_1__1__103_chanx_left_out;
wire [0:228] cbx_1__1__103_chanx_right_out;
wire [0:228] cbx_1__1__104_chanx_left_out;
wire [0:228] cbx_1__1__104_chanx_right_out;
wire [0:228] cbx_1__1__105_chanx_left_out;
wire [0:228] cbx_1__1__105_chanx_right_out;
wire [0:228] cbx_1__1__106_chanx_left_out;
wire [0:228] cbx_1__1__106_chanx_right_out;
wire [0:228] cbx_1__1__107_chanx_left_out;
wire [0:228] cbx_1__1__107_chanx_right_out;
wire [0:228] cbx_1__1__108_chanx_left_out;
wire [0:228] cbx_1__1__108_chanx_right_out;
wire [0:228] cbx_1__1__109_chanx_left_out;
wire [0:228] cbx_1__1__109_chanx_right_out;
wire [0:228] cbx_1__1__10_chanx_left_out;
wire [0:228] cbx_1__1__10_chanx_right_out;
wire [0:228] cbx_1__1__110_chanx_left_out;
wire [0:228] cbx_1__1__110_chanx_right_out;
wire [0:228] cbx_1__1__111_chanx_left_out;
wire [0:228] cbx_1__1__111_chanx_right_out;
wire [0:228] cbx_1__1__112_chanx_left_out;
wire [0:228] cbx_1__1__112_chanx_right_out;
wire [0:228] cbx_1__1__113_chanx_left_out;
wire [0:228] cbx_1__1__113_chanx_right_out;
wire [0:228] cbx_1__1__114_chanx_left_out;
wire [0:228] cbx_1__1__114_chanx_right_out;
wire [0:228] cbx_1__1__115_chanx_left_out;
wire [0:228] cbx_1__1__115_chanx_right_out;
wire [0:228] cbx_1__1__116_chanx_left_out;
wire [0:228] cbx_1__1__116_chanx_right_out;
wire [0:228] cbx_1__1__117_chanx_left_out;
wire [0:228] cbx_1__1__117_chanx_right_out;
wire [0:228] cbx_1__1__118_chanx_left_out;
wire [0:228] cbx_1__1__118_chanx_right_out;
wire [0:228] cbx_1__1__119_chanx_left_out;
wire [0:228] cbx_1__1__119_chanx_right_out;
wire [0:228] cbx_1__1__11_chanx_left_out;
wire [0:228] cbx_1__1__11_chanx_right_out;
wire [0:228] cbx_1__1__120_chanx_left_out;
wire [0:228] cbx_1__1__120_chanx_right_out;
wire [0:228] cbx_1__1__121_chanx_left_out;
wire [0:228] cbx_1__1__121_chanx_right_out;
wire [0:228] cbx_1__1__122_chanx_left_out;
wire [0:228] cbx_1__1__122_chanx_right_out;
wire [0:228] cbx_1__1__123_chanx_left_out;
wire [0:228] cbx_1__1__123_chanx_right_out;
wire [0:228] cbx_1__1__124_chanx_left_out;
wire [0:228] cbx_1__1__124_chanx_right_out;
wire [0:228] cbx_1__1__125_chanx_left_out;
wire [0:228] cbx_1__1__125_chanx_right_out;
wire [0:228] cbx_1__1__126_chanx_left_out;
wire [0:228] cbx_1__1__126_chanx_right_out;
wire [0:228] cbx_1__1__127_chanx_left_out;
wire [0:228] cbx_1__1__127_chanx_right_out;
wire [0:228] cbx_1__1__128_chanx_left_out;
wire [0:228] cbx_1__1__128_chanx_right_out;
wire [0:228] cbx_1__1__129_chanx_left_out;
wire [0:228] cbx_1__1__129_chanx_right_out;
wire [0:228] cbx_1__1__12_chanx_left_out;
wire [0:228] cbx_1__1__12_chanx_right_out;
wire [0:228] cbx_1__1__130_chanx_left_out;
wire [0:228] cbx_1__1__130_chanx_right_out;
wire [0:228] cbx_1__1__131_chanx_left_out;
wire [0:228] cbx_1__1__131_chanx_right_out;
wire [0:228] cbx_1__1__132_chanx_left_out;
wire [0:228] cbx_1__1__132_chanx_right_out;
wire [0:228] cbx_1__1__133_chanx_left_out;
wire [0:228] cbx_1__1__133_chanx_right_out;
wire [0:228] cbx_1__1__134_chanx_left_out;
wire [0:228] cbx_1__1__134_chanx_right_out;
wire [0:228] cbx_1__1__135_chanx_left_out;
wire [0:228] cbx_1__1__135_chanx_right_out;
wire [0:228] cbx_1__1__136_chanx_left_out;
wire [0:228] cbx_1__1__136_chanx_right_out;
wire [0:228] cbx_1__1__137_chanx_left_out;
wire [0:228] cbx_1__1__137_chanx_right_out;
wire [0:228] cbx_1__1__138_chanx_left_out;
wire [0:228] cbx_1__1__138_chanx_right_out;
wire [0:228] cbx_1__1__139_chanx_left_out;
wire [0:228] cbx_1__1__139_chanx_right_out;
wire [0:228] cbx_1__1__13_chanx_left_out;
wire [0:228] cbx_1__1__13_chanx_right_out;
wire [0:228] cbx_1__1__140_chanx_left_out;
wire [0:228] cbx_1__1__140_chanx_right_out;
wire [0:228] cbx_1__1__141_chanx_left_out;
wire [0:228] cbx_1__1__141_chanx_right_out;
wire [0:228] cbx_1__1__142_chanx_left_out;
wire [0:228] cbx_1__1__142_chanx_right_out;
wire [0:228] cbx_1__1__143_chanx_left_out;
wire [0:228] cbx_1__1__143_chanx_right_out;
wire [0:228] cbx_1__1__144_chanx_left_out;
wire [0:228] cbx_1__1__144_chanx_right_out;
wire [0:228] cbx_1__1__145_chanx_left_out;
wire [0:228] cbx_1__1__145_chanx_right_out;
wire [0:228] cbx_1__1__146_chanx_left_out;
wire [0:228] cbx_1__1__146_chanx_right_out;
wire [0:228] cbx_1__1__147_chanx_left_out;
wire [0:228] cbx_1__1__147_chanx_right_out;
wire [0:228] cbx_1__1__148_chanx_left_out;
wire [0:228] cbx_1__1__148_chanx_right_out;
wire [0:228] cbx_1__1__149_chanx_left_out;
wire [0:228] cbx_1__1__149_chanx_right_out;
wire [0:228] cbx_1__1__14_chanx_left_out;
wire [0:228] cbx_1__1__14_chanx_right_out;
wire [0:228] cbx_1__1__150_chanx_left_out;
wire [0:228] cbx_1__1__150_chanx_right_out;
wire [0:228] cbx_1__1__151_chanx_left_out;
wire [0:228] cbx_1__1__151_chanx_right_out;
wire [0:228] cbx_1__1__152_chanx_left_out;
wire [0:228] cbx_1__1__152_chanx_right_out;
wire [0:228] cbx_1__1__153_chanx_left_out;
wire [0:228] cbx_1__1__153_chanx_right_out;
wire [0:228] cbx_1__1__154_chanx_left_out;
wire [0:228] cbx_1__1__154_chanx_right_out;
wire [0:228] cbx_1__1__155_chanx_left_out;
wire [0:228] cbx_1__1__155_chanx_right_out;
wire [0:228] cbx_1__1__156_chanx_left_out;
wire [0:228] cbx_1__1__156_chanx_right_out;
wire [0:228] cbx_1__1__157_chanx_left_out;
wire [0:228] cbx_1__1__157_chanx_right_out;
wire [0:228] cbx_1__1__158_chanx_left_out;
wire [0:228] cbx_1__1__158_chanx_right_out;
wire [0:228] cbx_1__1__159_chanx_left_out;
wire [0:228] cbx_1__1__159_chanx_right_out;
wire [0:228] cbx_1__1__15_chanx_left_out;
wire [0:228] cbx_1__1__15_chanx_right_out;
wire [0:228] cbx_1__1__160_chanx_left_out;
wire [0:228] cbx_1__1__160_chanx_right_out;
wire [0:228] cbx_1__1__161_chanx_left_out;
wire [0:228] cbx_1__1__161_chanx_right_out;
wire [0:228] cbx_1__1__162_chanx_left_out;
wire [0:228] cbx_1__1__162_chanx_right_out;
wire [0:228] cbx_1__1__163_chanx_left_out;
wire [0:228] cbx_1__1__163_chanx_right_out;
wire [0:228] cbx_1__1__164_chanx_left_out;
wire [0:228] cbx_1__1__164_chanx_right_out;
wire [0:228] cbx_1__1__165_chanx_left_out;
wire [0:228] cbx_1__1__165_chanx_right_out;
wire [0:228] cbx_1__1__166_chanx_left_out;
wire [0:228] cbx_1__1__166_chanx_right_out;
wire [0:228] cbx_1__1__167_chanx_left_out;
wire [0:228] cbx_1__1__167_chanx_right_out;
wire [0:228] cbx_1__1__168_chanx_left_out;
wire [0:228] cbx_1__1__168_chanx_right_out;
wire [0:228] cbx_1__1__169_chanx_left_out;
wire [0:228] cbx_1__1__169_chanx_right_out;
wire [0:228] cbx_1__1__16_chanx_left_out;
wire [0:228] cbx_1__1__16_chanx_right_out;
wire [0:228] cbx_1__1__170_chanx_left_out;
wire [0:228] cbx_1__1__170_chanx_right_out;
wire [0:228] cbx_1__1__171_chanx_left_out;
wire [0:228] cbx_1__1__171_chanx_right_out;
wire [0:228] cbx_1__1__172_chanx_left_out;
wire [0:228] cbx_1__1__172_chanx_right_out;
wire [0:228] cbx_1__1__173_chanx_left_out;
wire [0:228] cbx_1__1__173_chanx_right_out;
wire [0:228] cbx_1__1__174_chanx_left_out;
wire [0:228] cbx_1__1__174_chanx_right_out;
wire [0:228] cbx_1__1__175_chanx_left_out;
wire [0:228] cbx_1__1__175_chanx_right_out;
wire [0:228] cbx_1__1__176_chanx_left_out;
wire [0:228] cbx_1__1__176_chanx_right_out;
wire [0:228] cbx_1__1__177_chanx_left_out;
wire [0:228] cbx_1__1__177_chanx_right_out;
wire [0:228] cbx_1__1__178_chanx_left_out;
wire [0:228] cbx_1__1__178_chanx_right_out;
wire [0:228] cbx_1__1__179_chanx_left_out;
wire [0:228] cbx_1__1__179_chanx_right_out;
wire [0:228] cbx_1__1__17_chanx_left_out;
wire [0:228] cbx_1__1__17_chanx_right_out;
wire [0:228] cbx_1__1__180_chanx_left_out;
wire [0:228] cbx_1__1__180_chanx_right_out;
wire [0:228] cbx_1__1__181_chanx_left_out;
wire [0:228] cbx_1__1__181_chanx_right_out;
wire [0:228] cbx_1__1__182_chanx_left_out;
wire [0:228] cbx_1__1__182_chanx_right_out;
wire [0:228] cbx_1__1__183_chanx_left_out;
wire [0:228] cbx_1__1__183_chanx_right_out;
wire [0:228] cbx_1__1__184_chanx_left_out;
wire [0:228] cbx_1__1__184_chanx_right_out;
wire [0:228] cbx_1__1__185_chanx_left_out;
wire [0:228] cbx_1__1__185_chanx_right_out;
wire [0:228] cbx_1__1__186_chanx_left_out;
wire [0:228] cbx_1__1__186_chanx_right_out;
wire [0:228] cbx_1__1__187_chanx_left_out;
wire [0:228] cbx_1__1__187_chanx_right_out;
wire [0:228] cbx_1__1__188_chanx_left_out;
wire [0:228] cbx_1__1__188_chanx_right_out;
wire [0:228] cbx_1__1__189_chanx_left_out;
wire [0:228] cbx_1__1__189_chanx_right_out;
wire [0:228] cbx_1__1__18_chanx_left_out;
wire [0:228] cbx_1__1__18_chanx_right_out;
wire [0:228] cbx_1__1__190_chanx_left_out;
wire [0:228] cbx_1__1__190_chanx_right_out;
wire [0:228] cbx_1__1__191_chanx_left_out;
wire [0:228] cbx_1__1__191_chanx_right_out;
wire [0:228] cbx_1__1__192_chanx_left_out;
wire [0:228] cbx_1__1__192_chanx_right_out;
wire [0:228] cbx_1__1__193_chanx_left_out;
wire [0:228] cbx_1__1__193_chanx_right_out;
wire [0:228] cbx_1__1__194_chanx_left_out;
wire [0:228] cbx_1__1__194_chanx_right_out;
wire [0:228] cbx_1__1__195_chanx_left_out;
wire [0:228] cbx_1__1__195_chanx_right_out;
wire [0:228] cbx_1__1__196_chanx_left_out;
wire [0:228] cbx_1__1__196_chanx_right_out;
wire [0:228] cbx_1__1__197_chanx_left_out;
wire [0:228] cbx_1__1__197_chanx_right_out;
wire [0:228] cbx_1__1__198_chanx_left_out;
wire [0:228] cbx_1__1__198_chanx_right_out;
wire [0:228] cbx_1__1__199_chanx_left_out;
wire [0:228] cbx_1__1__199_chanx_right_out;
wire [0:228] cbx_1__1__19_chanx_left_out;
wire [0:228] cbx_1__1__19_chanx_right_out;
wire [0:228] cbx_1__1__1_chanx_left_out;
wire [0:228] cbx_1__1__1_chanx_right_out;
wire [0:228] cbx_1__1__200_chanx_left_out;
wire [0:228] cbx_1__1__200_chanx_right_out;
wire [0:228] cbx_1__1__201_chanx_left_out;
wire [0:228] cbx_1__1__201_chanx_right_out;
wire [0:228] cbx_1__1__202_chanx_left_out;
wire [0:228] cbx_1__1__202_chanx_right_out;
wire [0:228] cbx_1__1__203_chanx_left_out;
wire [0:228] cbx_1__1__203_chanx_right_out;
wire [0:228] cbx_1__1__204_chanx_left_out;
wire [0:228] cbx_1__1__204_chanx_right_out;
wire [0:228] cbx_1__1__205_chanx_left_out;
wire [0:228] cbx_1__1__205_chanx_right_out;
wire [0:228] cbx_1__1__206_chanx_left_out;
wire [0:228] cbx_1__1__206_chanx_right_out;
wire [0:228] cbx_1__1__207_chanx_left_out;
wire [0:228] cbx_1__1__207_chanx_right_out;
wire [0:228] cbx_1__1__208_chanx_left_out;
wire [0:228] cbx_1__1__208_chanx_right_out;
wire [0:228] cbx_1__1__209_chanx_left_out;
wire [0:228] cbx_1__1__209_chanx_right_out;
wire [0:228] cbx_1__1__20_chanx_left_out;
wire [0:228] cbx_1__1__20_chanx_right_out;
wire [0:228] cbx_1__1__210_chanx_left_out;
wire [0:228] cbx_1__1__210_chanx_right_out;
wire [0:228] cbx_1__1__211_chanx_left_out;
wire [0:228] cbx_1__1__211_chanx_right_out;
wire [0:228] cbx_1__1__212_chanx_left_out;
wire [0:228] cbx_1__1__212_chanx_right_out;
wire [0:228] cbx_1__1__213_chanx_left_out;
wire [0:228] cbx_1__1__213_chanx_right_out;
wire [0:228] cbx_1__1__214_chanx_left_out;
wire [0:228] cbx_1__1__214_chanx_right_out;
wire [0:228] cbx_1__1__215_chanx_left_out;
wire [0:228] cbx_1__1__215_chanx_right_out;
wire [0:228] cbx_1__1__216_chanx_left_out;
wire [0:228] cbx_1__1__216_chanx_right_out;
wire [0:228] cbx_1__1__217_chanx_left_out;
wire [0:228] cbx_1__1__217_chanx_right_out;
wire [0:228] cbx_1__1__218_chanx_left_out;
wire [0:228] cbx_1__1__218_chanx_right_out;
wire [0:228] cbx_1__1__219_chanx_left_out;
wire [0:228] cbx_1__1__219_chanx_right_out;
wire [0:228] cbx_1__1__21_chanx_left_out;
wire [0:228] cbx_1__1__21_chanx_right_out;
wire [0:228] cbx_1__1__220_chanx_left_out;
wire [0:228] cbx_1__1__220_chanx_right_out;
wire [0:228] cbx_1__1__221_chanx_left_out;
wire [0:228] cbx_1__1__221_chanx_right_out;
wire [0:228] cbx_1__1__222_chanx_left_out;
wire [0:228] cbx_1__1__222_chanx_right_out;
wire [0:228] cbx_1__1__223_chanx_left_out;
wire [0:228] cbx_1__1__223_chanx_right_out;
wire [0:228] cbx_1__1__224_chanx_left_out;
wire [0:228] cbx_1__1__224_chanx_right_out;
wire [0:228] cbx_1__1__225_chanx_left_out;
wire [0:228] cbx_1__1__225_chanx_right_out;
wire [0:228] cbx_1__1__226_chanx_left_out;
wire [0:228] cbx_1__1__226_chanx_right_out;
wire [0:228] cbx_1__1__227_chanx_left_out;
wire [0:228] cbx_1__1__227_chanx_right_out;
wire [0:228] cbx_1__1__228_chanx_left_out;
wire [0:228] cbx_1__1__228_chanx_right_out;
wire [0:228] cbx_1__1__229_chanx_left_out;
wire [0:228] cbx_1__1__229_chanx_right_out;
wire [0:228] cbx_1__1__22_chanx_left_out;
wire [0:228] cbx_1__1__22_chanx_right_out;
wire [0:228] cbx_1__1__230_chanx_left_out;
wire [0:228] cbx_1__1__230_chanx_right_out;
wire [0:228] cbx_1__1__231_chanx_left_out;
wire [0:228] cbx_1__1__231_chanx_right_out;
wire [0:228] cbx_1__1__232_chanx_left_out;
wire [0:228] cbx_1__1__232_chanx_right_out;
wire [0:228] cbx_1__1__233_chanx_left_out;
wire [0:228] cbx_1__1__233_chanx_right_out;
wire [0:228] cbx_1__1__234_chanx_left_out;
wire [0:228] cbx_1__1__234_chanx_right_out;
wire [0:228] cbx_1__1__235_chanx_left_out;
wire [0:228] cbx_1__1__235_chanx_right_out;
wire [0:228] cbx_1__1__236_chanx_left_out;
wire [0:228] cbx_1__1__236_chanx_right_out;
wire [0:228] cbx_1__1__237_chanx_left_out;
wire [0:228] cbx_1__1__237_chanx_right_out;
wire [0:228] cbx_1__1__238_chanx_left_out;
wire [0:228] cbx_1__1__238_chanx_right_out;
wire [0:228] cbx_1__1__239_chanx_left_out;
wire [0:228] cbx_1__1__239_chanx_right_out;
wire [0:228] cbx_1__1__23_chanx_left_out;
wire [0:228] cbx_1__1__23_chanx_right_out;
wire [0:228] cbx_1__1__240_chanx_left_out;
wire [0:228] cbx_1__1__240_chanx_right_out;
wire [0:228] cbx_1__1__241_chanx_left_out;
wire [0:228] cbx_1__1__241_chanx_right_out;
wire [0:228] cbx_1__1__242_chanx_left_out;
wire [0:228] cbx_1__1__242_chanx_right_out;
wire [0:228] cbx_1__1__243_chanx_left_out;
wire [0:228] cbx_1__1__243_chanx_right_out;
wire [0:228] cbx_1__1__244_chanx_left_out;
wire [0:228] cbx_1__1__244_chanx_right_out;
wire [0:228] cbx_1__1__245_chanx_left_out;
wire [0:228] cbx_1__1__245_chanx_right_out;
wire [0:228] cbx_1__1__246_chanx_left_out;
wire [0:228] cbx_1__1__246_chanx_right_out;
wire [0:228] cbx_1__1__247_chanx_left_out;
wire [0:228] cbx_1__1__247_chanx_right_out;
wire [0:228] cbx_1__1__248_chanx_left_out;
wire [0:228] cbx_1__1__248_chanx_right_out;
wire [0:228] cbx_1__1__249_chanx_left_out;
wire [0:228] cbx_1__1__249_chanx_right_out;
wire [0:228] cbx_1__1__24_chanx_left_out;
wire [0:228] cbx_1__1__24_chanx_right_out;
wire [0:228] cbx_1__1__250_chanx_left_out;
wire [0:228] cbx_1__1__250_chanx_right_out;
wire [0:228] cbx_1__1__251_chanx_left_out;
wire [0:228] cbx_1__1__251_chanx_right_out;
wire [0:228] cbx_1__1__252_chanx_left_out;
wire [0:228] cbx_1__1__252_chanx_right_out;
wire [0:228] cbx_1__1__253_chanx_left_out;
wire [0:228] cbx_1__1__253_chanx_right_out;
wire [0:228] cbx_1__1__254_chanx_left_out;
wire [0:228] cbx_1__1__254_chanx_right_out;
wire [0:228] cbx_1__1__255_chanx_left_out;
wire [0:228] cbx_1__1__255_chanx_right_out;
wire [0:228] cbx_1__1__256_chanx_left_out;
wire [0:228] cbx_1__1__256_chanx_right_out;
wire [0:228] cbx_1__1__257_chanx_left_out;
wire [0:228] cbx_1__1__257_chanx_right_out;
wire [0:228] cbx_1__1__258_chanx_left_out;
wire [0:228] cbx_1__1__258_chanx_right_out;
wire [0:228] cbx_1__1__259_chanx_left_out;
wire [0:228] cbx_1__1__259_chanx_right_out;
wire [0:228] cbx_1__1__25_chanx_left_out;
wire [0:228] cbx_1__1__25_chanx_right_out;
wire [0:228] cbx_1__1__260_chanx_left_out;
wire [0:228] cbx_1__1__260_chanx_right_out;
wire [0:228] cbx_1__1__261_chanx_left_out;
wire [0:228] cbx_1__1__261_chanx_right_out;
wire [0:228] cbx_1__1__262_chanx_left_out;
wire [0:228] cbx_1__1__262_chanx_right_out;
wire [0:228] cbx_1__1__263_chanx_left_out;
wire [0:228] cbx_1__1__263_chanx_right_out;
wire [0:228] cbx_1__1__264_chanx_left_out;
wire [0:228] cbx_1__1__264_chanx_right_out;
wire [0:228] cbx_1__1__265_chanx_left_out;
wire [0:228] cbx_1__1__265_chanx_right_out;
wire [0:228] cbx_1__1__266_chanx_left_out;
wire [0:228] cbx_1__1__266_chanx_right_out;
wire [0:228] cbx_1__1__267_chanx_left_out;
wire [0:228] cbx_1__1__267_chanx_right_out;
wire [0:228] cbx_1__1__268_chanx_left_out;
wire [0:228] cbx_1__1__268_chanx_right_out;
wire [0:228] cbx_1__1__269_chanx_left_out;
wire [0:228] cbx_1__1__269_chanx_right_out;
wire [0:228] cbx_1__1__26_chanx_left_out;
wire [0:228] cbx_1__1__26_chanx_right_out;
wire [0:228] cbx_1__1__270_chanx_left_out;
wire [0:228] cbx_1__1__270_chanx_right_out;
wire [0:228] cbx_1__1__271_chanx_left_out;
wire [0:228] cbx_1__1__271_chanx_right_out;
wire [0:228] cbx_1__1__272_chanx_left_out;
wire [0:228] cbx_1__1__272_chanx_right_out;
wire [0:228] cbx_1__1__273_chanx_left_out;
wire [0:228] cbx_1__1__273_chanx_right_out;
wire [0:228] cbx_1__1__274_chanx_left_out;
wire [0:228] cbx_1__1__274_chanx_right_out;
wire [0:228] cbx_1__1__275_chanx_left_out;
wire [0:228] cbx_1__1__275_chanx_right_out;
wire [0:228] cbx_1__1__276_chanx_left_out;
wire [0:228] cbx_1__1__276_chanx_right_out;
wire [0:228] cbx_1__1__277_chanx_left_out;
wire [0:228] cbx_1__1__277_chanx_right_out;
wire [0:228] cbx_1__1__278_chanx_left_out;
wire [0:228] cbx_1__1__278_chanx_right_out;
wire [0:228] cbx_1__1__279_chanx_left_out;
wire [0:228] cbx_1__1__279_chanx_right_out;
wire [0:228] cbx_1__1__27_chanx_left_out;
wire [0:228] cbx_1__1__27_chanx_right_out;
wire [0:228] cbx_1__1__280_chanx_left_out;
wire [0:228] cbx_1__1__280_chanx_right_out;
wire [0:228] cbx_1__1__281_chanx_left_out;
wire [0:228] cbx_1__1__281_chanx_right_out;
wire [0:228] cbx_1__1__282_chanx_left_out;
wire [0:228] cbx_1__1__282_chanx_right_out;
wire [0:228] cbx_1__1__283_chanx_left_out;
wire [0:228] cbx_1__1__283_chanx_right_out;
wire [0:228] cbx_1__1__284_chanx_left_out;
wire [0:228] cbx_1__1__284_chanx_right_out;
wire [0:228] cbx_1__1__285_chanx_left_out;
wire [0:228] cbx_1__1__285_chanx_right_out;
wire [0:228] cbx_1__1__286_chanx_left_out;
wire [0:228] cbx_1__1__286_chanx_right_out;
wire [0:228] cbx_1__1__287_chanx_left_out;
wire [0:228] cbx_1__1__287_chanx_right_out;
wire [0:228] cbx_1__1__288_chanx_left_out;
wire [0:228] cbx_1__1__288_chanx_right_out;
wire [0:228] cbx_1__1__289_chanx_left_out;
wire [0:228] cbx_1__1__289_chanx_right_out;
wire [0:228] cbx_1__1__28_chanx_left_out;
wire [0:228] cbx_1__1__28_chanx_right_out;
wire [0:228] cbx_1__1__290_chanx_left_out;
wire [0:228] cbx_1__1__290_chanx_right_out;
wire [0:228] cbx_1__1__291_chanx_left_out;
wire [0:228] cbx_1__1__291_chanx_right_out;
wire [0:228] cbx_1__1__292_chanx_left_out;
wire [0:228] cbx_1__1__292_chanx_right_out;
wire [0:228] cbx_1__1__293_chanx_left_out;
wire [0:228] cbx_1__1__293_chanx_right_out;
wire [0:228] cbx_1__1__294_chanx_left_out;
wire [0:228] cbx_1__1__294_chanx_right_out;
wire [0:228] cbx_1__1__295_chanx_left_out;
wire [0:228] cbx_1__1__295_chanx_right_out;
wire [0:228] cbx_1__1__296_chanx_left_out;
wire [0:228] cbx_1__1__296_chanx_right_out;
wire [0:228] cbx_1__1__297_chanx_left_out;
wire [0:228] cbx_1__1__297_chanx_right_out;
wire [0:228] cbx_1__1__298_chanx_left_out;
wire [0:228] cbx_1__1__298_chanx_right_out;
wire [0:228] cbx_1__1__299_chanx_left_out;
wire [0:228] cbx_1__1__299_chanx_right_out;
wire [0:228] cbx_1__1__29_chanx_left_out;
wire [0:228] cbx_1__1__29_chanx_right_out;
wire [0:228] cbx_1__1__2_chanx_left_out;
wire [0:228] cbx_1__1__2_chanx_right_out;
wire [0:228] cbx_1__1__300_chanx_left_out;
wire [0:228] cbx_1__1__300_chanx_right_out;
wire [0:228] cbx_1__1__301_chanx_left_out;
wire [0:228] cbx_1__1__301_chanx_right_out;
wire [0:228] cbx_1__1__302_chanx_left_out;
wire [0:228] cbx_1__1__302_chanx_right_out;
wire [0:228] cbx_1__1__303_chanx_left_out;
wire [0:228] cbx_1__1__303_chanx_right_out;
wire [0:228] cbx_1__1__304_chanx_left_out;
wire [0:228] cbx_1__1__304_chanx_right_out;
wire [0:228] cbx_1__1__305_chanx_left_out;
wire [0:228] cbx_1__1__305_chanx_right_out;
wire [0:228] cbx_1__1__306_chanx_left_out;
wire [0:228] cbx_1__1__306_chanx_right_out;
wire [0:228] cbx_1__1__307_chanx_left_out;
wire [0:228] cbx_1__1__307_chanx_right_out;
wire [0:228] cbx_1__1__308_chanx_left_out;
wire [0:228] cbx_1__1__308_chanx_right_out;
wire [0:228] cbx_1__1__309_chanx_left_out;
wire [0:228] cbx_1__1__309_chanx_right_out;
wire [0:228] cbx_1__1__30_chanx_left_out;
wire [0:228] cbx_1__1__30_chanx_right_out;
wire [0:228] cbx_1__1__310_chanx_left_out;
wire [0:228] cbx_1__1__310_chanx_right_out;
wire [0:228] cbx_1__1__311_chanx_left_out;
wire [0:228] cbx_1__1__311_chanx_right_out;
wire [0:228] cbx_1__1__312_chanx_left_out;
wire [0:228] cbx_1__1__312_chanx_right_out;
wire [0:228] cbx_1__1__313_chanx_left_out;
wire [0:228] cbx_1__1__313_chanx_right_out;
wire [0:228] cbx_1__1__314_chanx_left_out;
wire [0:228] cbx_1__1__314_chanx_right_out;
wire [0:228] cbx_1__1__315_chanx_left_out;
wire [0:228] cbx_1__1__315_chanx_right_out;
wire [0:228] cbx_1__1__316_chanx_left_out;
wire [0:228] cbx_1__1__316_chanx_right_out;
wire [0:228] cbx_1__1__317_chanx_left_out;
wire [0:228] cbx_1__1__317_chanx_right_out;
wire [0:228] cbx_1__1__318_chanx_left_out;
wire [0:228] cbx_1__1__318_chanx_right_out;
wire [0:228] cbx_1__1__319_chanx_left_out;
wire [0:228] cbx_1__1__319_chanx_right_out;
wire [0:228] cbx_1__1__31_chanx_left_out;
wire [0:228] cbx_1__1__31_chanx_right_out;
wire [0:228] cbx_1__1__320_chanx_left_out;
wire [0:228] cbx_1__1__320_chanx_right_out;
wire [0:228] cbx_1__1__321_chanx_left_out;
wire [0:228] cbx_1__1__321_chanx_right_out;
wire [0:228] cbx_1__1__322_chanx_left_out;
wire [0:228] cbx_1__1__322_chanx_right_out;
wire [0:228] cbx_1__1__323_chanx_left_out;
wire [0:228] cbx_1__1__323_chanx_right_out;
wire [0:228] cbx_1__1__324_chanx_left_out;
wire [0:228] cbx_1__1__324_chanx_right_out;
wire [0:228] cbx_1__1__325_chanx_left_out;
wire [0:228] cbx_1__1__325_chanx_right_out;
wire [0:228] cbx_1__1__326_chanx_left_out;
wire [0:228] cbx_1__1__326_chanx_right_out;
wire [0:228] cbx_1__1__327_chanx_left_out;
wire [0:228] cbx_1__1__327_chanx_right_out;
wire [0:228] cbx_1__1__328_chanx_left_out;
wire [0:228] cbx_1__1__328_chanx_right_out;
wire [0:228] cbx_1__1__329_chanx_left_out;
wire [0:228] cbx_1__1__329_chanx_right_out;
wire [0:228] cbx_1__1__32_chanx_left_out;
wire [0:228] cbx_1__1__32_chanx_right_out;
wire [0:228] cbx_1__1__330_chanx_left_out;
wire [0:228] cbx_1__1__330_chanx_right_out;
wire [0:228] cbx_1__1__331_chanx_left_out;
wire [0:228] cbx_1__1__331_chanx_right_out;
wire [0:228] cbx_1__1__332_chanx_left_out;
wire [0:228] cbx_1__1__332_chanx_right_out;
wire [0:228] cbx_1__1__333_chanx_left_out;
wire [0:228] cbx_1__1__333_chanx_right_out;
wire [0:228] cbx_1__1__334_chanx_left_out;
wire [0:228] cbx_1__1__334_chanx_right_out;
wire [0:228] cbx_1__1__335_chanx_left_out;
wire [0:228] cbx_1__1__335_chanx_right_out;
wire [0:228] cbx_1__1__336_chanx_left_out;
wire [0:228] cbx_1__1__336_chanx_right_out;
wire [0:228] cbx_1__1__337_chanx_left_out;
wire [0:228] cbx_1__1__337_chanx_right_out;
wire [0:228] cbx_1__1__338_chanx_left_out;
wire [0:228] cbx_1__1__338_chanx_right_out;
wire [0:228] cbx_1__1__339_chanx_left_out;
wire [0:228] cbx_1__1__339_chanx_right_out;
wire [0:228] cbx_1__1__33_chanx_left_out;
wire [0:228] cbx_1__1__33_chanx_right_out;
wire [0:228] cbx_1__1__340_chanx_left_out;
wire [0:228] cbx_1__1__340_chanx_right_out;
wire [0:228] cbx_1__1__341_chanx_left_out;
wire [0:228] cbx_1__1__341_chanx_right_out;
wire [0:228] cbx_1__1__342_chanx_left_out;
wire [0:228] cbx_1__1__342_chanx_right_out;
wire [0:228] cbx_1__1__343_chanx_left_out;
wire [0:228] cbx_1__1__343_chanx_right_out;
wire [0:228] cbx_1__1__344_chanx_left_out;
wire [0:228] cbx_1__1__344_chanx_right_out;
wire [0:228] cbx_1__1__345_chanx_left_out;
wire [0:228] cbx_1__1__345_chanx_right_out;
wire [0:228] cbx_1__1__346_chanx_left_out;
wire [0:228] cbx_1__1__346_chanx_right_out;
wire [0:228] cbx_1__1__347_chanx_left_out;
wire [0:228] cbx_1__1__347_chanx_right_out;
wire [0:228] cbx_1__1__348_chanx_left_out;
wire [0:228] cbx_1__1__348_chanx_right_out;
wire [0:228] cbx_1__1__349_chanx_left_out;
wire [0:228] cbx_1__1__349_chanx_right_out;
wire [0:228] cbx_1__1__34_chanx_left_out;
wire [0:228] cbx_1__1__34_chanx_right_out;
wire [0:228] cbx_1__1__350_chanx_left_out;
wire [0:228] cbx_1__1__350_chanx_right_out;
wire [0:228] cbx_1__1__351_chanx_left_out;
wire [0:228] cbx_1__1__351_chanx_right_out;
wire [0:228] cbx_1__1__352_chanx_left_out;
wire [0:228] cbx_1__1__352_chanx_right_out;
wire [0:228] cbx_1__1__353_chanx_left_out;
wire [0:228] cbx_1__1__353_chanx_right_out;
wire [0:228] cbx_1__1__354_chanx_left_out;
wire [0:228] cbx_1__1__354_chanx_right_out;
wire [0:228] cbx_1__1__355_chanx_left_out;
wire [0:228] cbx_1__1__355_chanx_right_out;
wire [0:228] cbx_1__1__356_chanx_left_out;
wire [0:228] cbx_1__1__356_chanx_right_out;
wire [0:228] cbx_1__1__357_chanx_left_out;
wire [0:228] cbx_1__1__357_chanx_right_out;
wire [0:228] cbx_1__1__358_chanx_left_out;
wire [0:228] cbx_1__1__358_chanx_right_out;
wire [0:228] cbx_1__1__359_chanx_left_out;
wire [0:228] cbx_1__1__359_chanx_right_out;
wire [0:228] cbx_1__1__35_chanx_left_out;
wire [0:228] cbx_1__1__35_chanx_right_out;
wire [0:228] cbx_1__1__360_chanx_left_out;
wire [0:228] cbx_1__1__360_chanx_right_out;
wire [0:228] cbx_1__1__361_chanx_left_out;
wire [0:228] cbx_1__1__361_chanx_right_out;
wire [0:228] cbx_1__1__362_chanx_left_out;
wire [0:228] cbx_1__1__362_chanx_right_out;
wire [0:228] cbx_1__1__363_chanx_left_out;
wire [0:228] cbx_1__1__363_chanx_right_out;
wire [0:228] cbx_1__1__364_chanx_left_out;
wire [0:228] cbx_1__1__364_chanx_right_out;
wire [0:228] cbx_1__1__365_chanx_left_out;
wire [0:228] cbx_1__1__365_chanx_right_out;
wire [0:228] cbx_1__1__366_chanx_left_out;
wire [0:228] cbx_1__1__366_chanx_right_out;
wire [0:228] cbx_1__1__367_chanx_left_out;
wire [0:228] cbx_1__1__367_chanx_right_out;
wire [0:228] cbx_1__1__368_chanx_left_out;
wire [0:228] cbx_1__1__368_chanx_right_out;
wire [0:228] cbx_1__1__369_chanx_left_out;
wire [0:228] cbx_1__1__369_chanx_right_out;
wire [0:228] cbx_1__1__36_chanx_left_out;
wire [0:228] cbx_1__1__36_chanx_right_out;
wire [0:228] cbx_1__1__370_chanx_left_out;
wire [0:228] cbx_1__1__370_chanx_right_out;
wire [0:228] cbx_1__1__371_chanx_left_out;
wire [0:228] cbx_1__1__371_chanx_right_out;
wire [0:228] cbx_1__1__372_chanx_left_out;
wire [0:228] cbx_1__1__372_chanx_right_out;
wire [0:228] cbx_1__1__373_chanx_left_out;
wire [0:228] cbx_1__1__373_chanx_right_out;
wire [0:228] cbx_1__1__374_chanx_left_out;
wire [0:228] cbx_1__1__374_chanx_right_out;
wire [0:228] cbx_1__1__375_chanx_left_out;
wire [0:228] cbx_1__1__375_chanx_right_out;
wire [0:228] cbx_1__1__376_chanx_left_out;
wire [0:228] cbx_1__1__376_chanx_right_out;
wire [0:228] cbx_1__1__377_chanx_left_out;
wire [0:228] cbx_1__1__377_chanx_right_out;
wire [0:228] cbx_1__1__378_chanx_left_out;
wire [0:228] cbx_1__1__378_chanx_right_out;
wire [0:228] cbx_1__1__379_chanx_left_out;
wire [0:228] cbx_1__1__379_chanx_right_out;
wire [0:228] cbx_1__1__37_chanx_left_out;
wire [0:228] cbx_1__1__37_chanx_right_out;
wire [0:228] cbx_1__1__380_chanx_left_out;
wire [0:228] cbx_1__1__380_chanx_right_out;
wire [0:228] cbx_1__1__381_chanx_left_out;
wire [0:228] cbx_1__1__381_chanx_right_out;
wire [0:228] cbx_1__1__382_chanx_left_out;
wire [0:228] cbx_1__1__382_chanx_right_out;
wire [0:228] cbx_1__1__383_chanx_left_out;
wire [0:228] cbx_1__1__383_chanx_right_out;
wire [0:228] cbx_1__1__384_chanx_left_out;
wire [0:228] cbx_1__1__384_chanx_right_out;
wire [0:228] cbx_1__1__385_chanx_left_out;
wire [0:228] cbx_1__1__385_chanx_right_out;
wire [0:228] cbx_1__1__386_chanx_left_out;
wire [0:228] cbx_1__1__386_chanx_right_out;
wire [0:228] cbx_1__1__387_chanx_left_out;
wire [0:228] cbx_1__1__387_chanx_right_out;
wire [0:228] cbx_1__1__388_chanx_left_out;
wire [0:228] cbx_1__1__388_chanx_right_out;
wire [0:228] cbx_1__1__389_chanx_left_out;
wire [0:228] cbx_1__1__389_chanx_right_out;
wire [0:228] cbx_1__1__38_chanx_left_out;
wire [0:228] cbx_1__1__38_chanx_right_out;
wire [0:228] cbx_1__1__390_chanx_left_out;
wire [0:228] cbx_1__1__390_chanx_right_out;
wire [0:228] cbx_1__1__391_chanx_left_out;
wire [0:228] cbx_1__1__391_chanx_right_out;
wire [0:228] cbx_1__1__392_chanx_left_out;
wire [0:228] cbx_1__1__392_chanx_right_out;
wire [0:228] cbx_1__1__393_chanx_left_out;
wire [0:228] cbx_1__1__393_chanx_right_out;
wire [0:228] cbx_1__1__394_chanx_left_out;
wire [0:228] cbx_1__1__394_chanx_right_out;
wire [0:228] cbx_1__1__395_chanx_left_out;
wire [0:228] cbx_1__1__395_chanx_right_out;
wire [0:228] cbx_1__1__396_chanx_left_out;
wire [0:228] cbx_1__1__396_chanx_right_out;
wire [0:228] cbx_1__1__397_chanx_left_out;
wire [0:228] cbx_1__1__397_chanx_right_out;
wire [0:228] cbx_1__1__398_chanx_left_out;
wire [0:228] cbx_1__1__398_chanx_right_out;
wire [0:228] cbx_1__1__399_chanx_left_out;
wire [0:228] cbx_1__1__399_chanx_right_out;
wire [0:228] cbx_1__1__39_chanx_left_out;
wire [0:228] cbx_1__1__39_chanx_right_out;
wire [0:228] cbx_1__1__3_chanx_left_out;
wire [0:228] cbx_1__1__3_chanx_right_out;
wire [0:228] cbx_1__1__400_chanx_left_out;
wire [0:228] cbx_1__1__400_chanx_right_out;
wire [0:228] cbx_1__1__401_chanx_left_out;
wire [0:228] cbx_1__1__401_chanx_right_out;
wire [0:228] cbx_1__1__402_chanx_left_out;
wire [0:228] cbx_1__1__402_chanx_right_out;
wire [0:228] cbx_1__1__40_chanx_left_out;
wire [0:228] cbx_1__1__40_chanx_right_out;
wire [0:228] cbx_1__1__41_chanx_left_out;
wire [0:228] cbx_1__1__41_chanx_right_out;
wire [0:228] cbx_1__1__42_chanx_left_out;
wire [0:228] cbx_1__1__42_chanx_right_out;
wire [0:228] cbx_1__1__43_chanx_left_out;
wire [0:228] cbx_1__1__43_chanx_right_out;
wire [0:228] cbx_1__1__44_chanx_left_out;
wire [0:228] cbx_1__1__44_chanx_right_out;
wire [0:228] cbx_1__1__45_chanx_left_out;
wire [0:228] cbx_1__1__45_chanx_right_out;
wire [0:228] cbx_1__1__46_chanx_left_out;
wire [0:228] cbx_1__1__46_chanx_right_out;
wire [0:228] cbx_1__1__47_chanx_left_out;
wire [0:228] cbx_1__1__47_chanx_right_out;
wire [0:228] cbx_1__1__48_chanx_left_out;
wire [0:228] cbx_1__1__48_chanx_right_out;
wire [0:228] cbx_1__1__49_chanx_left_out;
wire [0:228] cbx_1__1__49_chanx_right_out;
wire [0:228] cbx_1__1__4_chanx_left_out;
wire [0:228] cbx_1__1__4_chanx_right_out;
wire [0:228] cbx_1__1__50_chanx_left_out;
wire [0:228] cbx_1__1__50_chanx_right_out;
wire [0:228] cbx_1__1__51_chanx_left_out;
wire [0:228] cbx_1__1__51_chanx_right_out;
wire [0:228] cbx_1__1__52_chanx_left_out;
wire [0:228] cbx_1__1__52_chanx_right_out;
wire [0:228] cbx_1__1__53_chanx_left_out;
wire [0:228] cbx_1__1__53_chanx_right_out;
wire [0:228] cbx_1__1__54_chanx_left_out;
wire [0:228] cbx_1__1__54_chanx_right_out;
wire [0:228] cbx_1__1__55_chanx_left_out;
wire [0:228] cbx_1__1__55_chanx_right_out;
wire [0:228] cbx_1__1__56_chanx_left_out;
wire [0:228] cbx_1__1__56_chanx_right_out;
wire [0:228] cbx_1__1__57_chanx_left_out;
wire [0:228] cbx_1__1__57_chanx_right_out;
wire [0:228] cbx_1__1__58_chanx_left_out;
wire [0:228] cbx_1__1__58_chanx_right_out;
wire [0:228] cbx_1__1__59_chanx_left_out;
wire [0:228] cbx_1__1__59_chanx_right_out;
wire [0:228] cbx_1__1__5_chanx_left_out;
wire [0:228] cbx_1__1__5_chanx_right_out;
wire [0:228] cbx_1__1__60_chanx_left_out;
wire [0:228] cbx_1__1__60_chanx_right_out;
wire [0:228] cbx_1__1__61_chanx_left_out;
wire [0:228] cbx_1__1__61_chanx_right_out;
wire [0:228] cbx_1__1__62_chanx_left_out;
wire [0:228] cbx_1__1__62_chanx_right_out;
wire [0:228] cbx_1__1__63_chanx_left_out;
wire [0:228] cbx_1__1__63_chanx_right_out;
wire [0:228] cbx_1__1__64_chanx_left_out;
wire [0:228] cbx_1__1__64_chanx_right_out;
wire [0:228] cbx_1__1__65_chanx_left_out;
wire [0:228] cbx_1__1__65_chanx_right_out;
wire [0:228] cbx_1__1__66_chanx_left_out;
wire [0:228] cbx_1__1__66_chanx_right_out;
wire [0:228] cbx_1__1__67_chanx_left_out;
wire [0:228] cbx_1__1__67_chanx_right_out;
wire [0:228] cbx_1__1__68_chanx_left_out;
wire [0:228] cbx_1__1__68_chanx_right_out;
wire [0:228] cbx_1__1__69_chanx_left_out;
wire [0:228] cbx_1__1__69_chanx_right_out;
wire [0:228] cbx_1__1__6_chanx_left_out;
wire [0:228] cbx_1__1__6_chanx_right_out;
wire [0:228] cbx_1__1__70_chanx_left_out;
wire [0:228] cbx_1__1__70_chanx_right_out;
wire [0:228] cbx_1__1__71_chanx_left_out;
wire [0:228] cbx_1__1__71_chanx_right_out;
wire [0:228] cbx_1__1__72_chanx_left_out;
wire [0:228] cbx_1__1__72_chanx_right_out;
wire [0:228] cbx_1__1__73_chanx_left_out;
wire [0:228] cbx_1__1__73_chanx_right_out;
wire [0:228] cbx_1__1__74_chanx_left_out;
wire [0:228] cbx_1__1__74_chanx_right_out;
wire [0:228] cbx_1__1__75_chanx_left_out;
wire [0:228] cbx_1__1__75_chanx_right_out;
wire [0:228] cbx_1__1__76_chanx_left_out;
wire [0:228] cbx_1__1__76_chanx_right_out;
wire [0:228] cbx_1__1__77_chanx_left_out;
wire [0:228] cbx_1__1__77_chanx_right_out;
wire [0:228] cbx_1__1__78_chanx_left_out;
wire [0:228] cbx_1__1__78_chanx_right_out;
wire [0:228] cbx_1__1__79_chanx_left_out;
wire [0:228] cbx_1__1__79_chanx_right_out;
wire [0:228] cbx_1__1__7_chanx_left_out;
wire [0:228] cbx_1__1__7_chanx_right_out;
wire [0:228] cbx_1__1__80_chanx_left_out;
wire [0:228] cbx_1__1__80_chanx_right_out;
wire [0:228] cbx_1__1__81_chanx_left_out;
wire [0:228] cbx_1__1__81_chanx_right_out;
wire [0:228] cbx_1__1__82_chanx_left_out;
wire [0:228] cbx_1__1__82_chanx_right_out;
wire [0:228] cbx_1__1__83_chanx_left_out;
wire [0:228] cbx_1__1__83_chanx_right_out;
wire [0:228] cbx_1__1__84_chanx_left_out;
wire [0:228] cbx_1__1__84_chanx_right_out;
wire [0:228] cbx_1__1__85_chanx_left_out;
wire [0:228] cbx_1__1__85_chanx_right_out;
wire [0:228] cbx_1__1__86_chanx_left_out;
wire [0:228] cbx_1__1__86_chanx_right_out;
wire [0:228] cbx_1__1__87_chanx_left_out;
wire [0:228] cbx_1__1__87_chanx_right_out;
wire [0:228] cbx_1__1__88_chanx_left_out;
wire [0:228] cbx_1__1__88_chanx_right_out;
wire [0:228] cbx_1__1__89_chanx_left_out;
wire [0:228] cbx_1__1__89_chanx_right_out;
wire [0:228] cbx_1__1__8_chanx_left_out;
wire [0:228] cbx_1__1__8_chanx_right_out;
wire [0:228] cbx_1__1__90_chanx_left_out;
wire [0:228] cbx_1__1__90_chanx_right_out;
wire [0:228] cbx_1__1__91_chanx_left_out;
wire [0:228] cbx_1__1__91_chanx_right_out;
wire [0:228] cbx_1__1__92_chanx_left_out;
wire [0:228] cbx_1__1__92_chanx_right_out;
wire [0:228] cbx_1__1__93_chanx_left_out;
wire [0:228] cbx_1__1__93_chanx_right_out;
wire [0:228] cbx_1__1__94_chanx_left_out;
wire [0:228] cbx_1__1__94_chanx_right_out;
wire [0:228] cbx_1__1__95_chanx_left_out;
wire [0:228] cbx_1__1__95_chanx_right_out;
wire [0:228] cbx_1__1__96_chanx_left_out;
wire [0:228] cbx_1__1__96_chanx_right_out;
wire [0:228] cbx_1__1__97_chanx_left_out;
wire [0:228] cbx_1__1__97_chanx_right_out;
wire [0:228] cbx_1__1__98_chanx_left_out;
wire [0:228] cbx_1__1__98_chanx_right_out;
wire [0:228] cbx_1__1__99_chanx_left_out;
wire [0:228] cbx_1__1__99_chanx_right_out;
wire [0:228] cbx_1__1__9_chanx_left_out;
wire [0:228] cbx_1__1__9_chanx_right_out;
wire [0:0] cbx_1__22__0_ccff_tail;
wire [0:228] cbx_1__22__0_chanx_left_out;
wire [0:228] cbx_1__22__0_chanx_right_out;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__10_ccff_tail;
wire [0:228] cbx_1__22__10_chanx_left_out;
wire [0:228] cbx_1__22__10_chanx_right_out;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__11_ccff_tail;
wire [0:228] cbx_1__22__11_chanx_left_out;
wire [0:228] cbx_1__22__11_chanx_right_out;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__12_ccff_tail;
wire [0:228] cbx_1__22__12_chanx_left_out;
wire [0:228] cbx_1__22__12_chanx_right_out;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__13_ccff_tail;
wire [0:228] cbx_1__22__13_chanx_left_out;
wire [0:228] cbx_1__22__13_chanx_right_out;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__14_ccff_tail;
wire [0:228] cbx_1__22__14_chanx_left_out;
wire [0:228] cbx_1__22__14_chanx_right_out;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__15_ccff_tail;
wire [0:228] cbx_1__22__15_chanx_left_out;
wire [0:228] cbx_1__22__15_chanx_right_out;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__16_ccff_tail;
wire [0:228] cbx_1__22__16_chanx_left_out;
wire [0:228] cbx_1__22__16_chanx_right_out;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__17_ccff_tail;
wire [0:228] cbx_1__22__17_chanx_left_out;
wire [0:228] cbx_1__22__17_chanx_right_out;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__18_ccff_tail;
wire [0:228] cbx_1__22__18_chanx_left_out;
wire [0:228] cbx_1__22__18_chanx_right_out;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__19_ccff_tail;
wire [0:228] cbx_1__22__19_chanx_left_out;
wire [0:228] cbx_1__22__19_chanx_right_out;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__1_ccff_tail;
wire [0:228] cbx_1__22__1_chanx_left_out;
wire [0:228] cbx_1__22__1_chanx_right_out;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__20_ccff_tail;
wire [0:228] cbx_1__22__20_chanx_left_out;
wire [0:228] cbx_1__22__20_chanx_right_out;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__21_ccff_tail;
wire [0:228] cbx_1__22__21_chanx_left_out;
wire [0:228] cbx_1__22__21_chanx_right_out;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__2_ccff_tail;
wire [0:228] cbx_1__22__2_chanx_left_out;
wire [0:228] cbx_1__22__2_chanx_right_out;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__3_ccff_tail;
wire [0:228] cbx_1__22__3_chanx_left_out;
wire [0:228] cbx_1__22__3_chanx_right_out;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__4_ccff_tail;
wire [0:228] cbx_1__22__4_chanx_left_out;
wire [0:228] cbx_1__22__4_chanx_right_out;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__5_ccff_tail;
wire [0:228] cbx_1__22__5_chanx_left_out;
wire [0:228] cbx_1__22__5_chanx_right_out;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__6_ccff_tail;
wire [0:228] cbx_1__22__6_chanx_left_out;
wire [0:228] cbx_1__22__6_chanx_right_out;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__7_ccff_tail;
wire [0:228] cbx_1__22__7_chanx_left_out;
wire [0:228] cbx_1__22__7_chanx_right_out;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__8_ccff_tail;
wire [0:228] cbx_1__22__8_chanx_left_out;
wire [0:228] cbx_1__22__8_chanx_right_out;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__22__9_ccff_tail;
wire [0:228] cbx_1__22__9_chanx_left_out;
wire [0:228] cbx_1__22__9_chanx_right_out;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__4__0_ccff_tail;
wire [0:228] cbx_1__4__0_chanx_left_out;
wire [0:228] cbx_1__4__0_chanx_right_out;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__10_ccff_tail;
wire [0:228] cbx_1__4__10_chanx_left_out;
wire [0:228] cbx_1__4__10_chanx_right_out;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__11_ccff_tail;
wire [0:228] cbx_1__4__11_chanx_left_out;
wire [0:228] cbx_1__4__11_chanx_right_out;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__12_ccff_tail;
wire [0:228] cbx_1__4__12_chanx_left_out;
wire [0:228] cbx_1__4__12_chanx_right_out;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__13_ccff_tail;
wire [0:228] cbx_1__4__13_chanx_left_out;
wire [0:228] cbx_1__4__13_chanx_right_out;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__14_ccff_tail;
wire [0:228] cbx_1__4__14_chanx_left_out;
wire [0:228] cbx_1__4__14_chanx_right_out;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__15_ccff_tail;
wire [0:228] cbx_1__4__15_chanx_left_out;
wire [0:228] cbx_1__4__15_chanx_right_out;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__16_ccff_tail;
wire [0:228] cbx_1__4__16_chanx_left_out;
wire [0:228] cbx_1__4__16_chanx_right_out;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__17_ccff_tail;
wire [0:228] cbx_1__4__17_chanx_left_out;
wire [0:228] cbx_1__4__17_chanx_right_out;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__18_ccff_tail;
wire [0:228] cbx_1__4__18_chanx_left_out;
wire [0:228] cbx_1__4__18_chanx_right_out;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__19_ccff_tail;
wire [0:228] cbx_1__4__19_chanx_left_out;
wire [0:228] cbx_1__4__19_chanx_right_out;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__1_ccff_tail;
wire [0:228] cbx_1__4__1_chanx_left_out;
wire [0:228] cbx_1__4__1_chanx_right_out;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__20_ccff_tail;
wire [0:228] cbx_1__4__20_chanx_left_out;
wire [0:228] cbx_1__4__20_chanx_right_out;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__21_ccff_tail;
wire [0:228] cbx_1__4__21_chanx_left_out;
wire [0:228] cbx_1__4__21_chanx_right_out;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__2_ccff_tail;
wire [0:228] cbx_1__4__2_chanx_left_out;
wire [0:228] cbx_1__4__2_chanx_right_out;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__3_ccff_tail;
wire [0:228] cbx_1__4__3_chanx_left_out;
wire [0:228] cbx_1__4__3_chanx_right_out;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__4_ccff_tail;
wire [0:228] cbx_1__4__4_chanx_left_out;
wire [0:228] cbx_1__4__4_chanx_right_out;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__5_ccff_tail;
wire [0:228] cbx_1__4__5_chanx_left_out;
wire [0:228] cbx_1__4__5_chanx_right_out;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__6_ccff_tail;
wire [0:228] cbx_1__4__6_chanx_left_out;
wire [0:228] cbx_1__4__6_chanx_right_out;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__7_ccff_tail;
wire [0:228] cbx_1__4__7_chanx_left_out;
wire [0:228] cbx_1__4__7_chanx_right_out;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__8_ccff_tail;
wire [0:228] cbx_1__4__8_chanx_left_out;
wire [0:228] cbx_1__4__8_chanx_right_out;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__4__9_ccff_tail;
wire [0:228] cbx_1__4__9_chanx_left_out;
wire [0:228] cbx_1__4__9_chanx_right_out;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__0_ccff_tail;
wire [0:228] cbx_1__5__0_chanx_left_out;
wire [0:228] cbx_1__5__0_chanx_right_out;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__10_ccff_tail;
wire [0:228] cbx_1__5__10_chanx_left_out;
wire [0:228] cbx_1__5__10_chanx_right_out;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__11_ccff_tail;
wire [0:228] cbx_1__5__11_chanx_left_out;
wire [0:228] cbx_1__5__11_chanx_right_out;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__12_ccff_tail;
wire [0:228] cbx_1__5__12_chanx_left_out;
wire [0:228] cbx_1__5__12_chanx_right_out;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__13_ccff_tail;
wire [0:228] cbx_1__5__13_chanx_left_out;
wire [0:228] cbx_1__5__13_chanx_right_out;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__14_ccff_tail;
wire [0:228] cbx_1__5__14_chanx_left_out;
wire [0:228] cbx_1__5__14_chanx_right_out;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__15_ccff_tail;
wire [0:228] cbx_1__5__15_chanx_left_out;
wire [0:228] cbx_1__5__15_chanx_right_out;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__16_ccff_tail;
wire [0:228] cbx_1__5__16_chanx_left_out;
wire [0:228] cbx_1__5__16_chanx_right_out;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__17_ccff_tail;
wire [0:228] cbx_1__5__17_chanx_left_out;
wire [0:228] cbx_1__5__17_chanx_right_out;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__18_ccff_tail;
wire [0:228] cbx_1__5__18_chanx_left_out;
wire [0:228] cbx_1__5__18_chanx_right_out;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__1_ccff_tail;
wire [0:228] cbx_1__5__1_chanx_left_out;
wire [0:228] cbx_1__5__1_chanx_right_out;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__2_ccff_tail;
wire [0:228] cbx_1__5__2_chanx_left_out;
wire [0:228] cbx_1__5__2_chanx_right_out;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__3_ccff_tail;
wire [0:228] cbx_1__5__3_chanx_left_out;
wire [0:228] cbx_1__5__3_chanx_right_out;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__4_ccff_tail;
wire [0:228] cbx_1__5__4_chanx_left_out;
wire [0:228] cbx_1__5__4_chanx_right_out;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__5_ccff_tail;
wire [0:228] cbx_1__5__5_chanx_left_out;
wire [0:228] cbx_1__5__5_chanx_right_out;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__6_ccff_tail;
wire [0:228] cbx_1__5__6_chanx_left_out;
wire [0:228] cbx_1__5__6_chanx_right_out;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__7_ccff_tail;
wire [0:228] cbx_1__5__7_chanx_left_out;
wire [0:228] cbx_1__5__7_chanx_right_out;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__8_ccff_tail;
wire [0:228] cbx_1__5__8_chanx_left_out;
wire [0:228] cbx_1__5__8_chanx_right_out;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__5__9_ccff_tail;
wire [0:228] cbx_1__5__9_chanx_left_out;
wire [0:228] cbx_1__5__9_chanx_right_out;
wire [0:0] cbx_3__2__0_ccff_tail;
wire [0:228] cbx_3__2__0_chanx_left_out;
wire [0:228] cbx_3__2__0_chanx_right_out;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__2__1_ccff_tail;
wire [0:228] cbx_3__2__1_chanx_left_out;
wire [0:228] cbx_3__2__1_chanx_right_out;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__2__2_ccff_tail;
wire [0:228] cbx_3__2__2_chanx_left_out;
wire [0:228] cbx_3__2__2_chanx_right_out;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__2__3_ccff_tail;
wire [0:228] cbx_3__2__3_chanx_left_out;
wire [0:228] cbx_3__2__3_chanx_right_out;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__2__4_ccff_tail;
wire [0:228] cbx_3__2__4_chanx_left_out;
wire [0:228] cbx_3__2__4_chanx_right_out;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__2__5_ccff_tail;
wire [0:228] cbx_3__2__5_chanx_left_out;
wire [0:228] cbx_3__2__5_chanx_right_out;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__0_ccff_tail;
wire [0:228] cbx_3__3__0_chanx_left_out;
wire [0:228] cbx_3__3__0_chanx_right_out;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__1_ccff_tail;
wire [0:228] cbx_3__3__1_chanx_left_out;
wire [0:228] cbx_3__3__1_chanx_right_out;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__2_ccff_tail;
wire [0:228] cbx_3__3__2_chanx_left_out;
wire [0:228] cbx_3__3__2_chanx_right_out;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__3_ccff_tail;
wire [0:228] cbx_3__3__3_chanx_left_out;
wire [0:228] cbx_3__3__3_chanx_right_out;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__4_ccff_tail;
wire [0:228] cbx_3__3__4_chanx_left_out;
wire [0:228] cbx_3__3__4_chanx_right_out;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__5_ccff_tail;
wire [0:228] cbx_3__3__5_chanx_left_out;
wire [0:228] cbx_3__3__5_chanx_right_out;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__6_ccff_tail;
wire [0:228] cbx_3__3__6_chanx_left_out;
wire [0:228] cbx_3__3__6_chanx_right_out;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__7_ccff_tail;
wire [0:228] cbx_3__3__7_chanx_left_out;
wire [0:228] cbx_3__3__7_chanx_right_out;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cbx_3__3__8_ccff_tail;
wire [0:228] cbx_3__3__8_chanx_left_out;
wire [0:228] cbx_3__3__8_chanx_right_out;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_3__5__0_ccff_tail;
wire [0:228] cbx_3__5__0_chanx_left_out;
wire [0:228] cbx_3__5__0_chanx_right_out;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_3__5__1_ccff_tail;
wire [0:228] cbx_3__5__1_chanx_left_out;
wire [0:228] cbx_3__5__1_chanx_right_out;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_3__5__2_ccff_tail;
wire [0:228] cbx_3__5__2_chanx_left_out;
wire [0:228] cbx_3__5__2_chanx_right_out;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:228] cby_0__1__0_chany_bottom_out;
wire [0:228] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__10_ccff_tail;
wire [0:228] cby_0__1__10_chany_bottom_out;
wire [0:228] cby_0__1__10_chany_top_out;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__11_ccff_tail;
wire [0:228] cby_0__1__11_chany_bottom_out;
wire [0:228] cby_0__1__11_chany_top_out;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__12_ccff_tail;
wire [0:228] cby_0__1__12_chany_bottom_out;
wire [0:228] cby_0__1__12_chany_top_out;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__13_ccff_tail;
wire [0:228] cby_0__1__13_chany_bottom_out;
wire [0:228] cby_0__1__13_chany_top_out;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__14_ccff_tail;
wire [0:228] cby_0__1__14_chany_bottom_out;
wire [0:228] cby_0__1__14_chany_top_out;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__15_ccff_tail;
wire [0:228] cby_0__1__15_chany_bottom_out;
wire [0:228] cby_0__1__15_chany_top_out;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__16_ccff_tail;
wire [0:228] cby_0__1__16_chany_bottom_out;
wire [0:228] cby_0__1__16_chany_top_out;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__17_ccff_tail;
wire [0:228] cby_0__1__17_chany_bottom_out;
wire [0:228] cby_0__1__17_chany_top_out;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__18_ccff_tail;
wire [0:228] cby_0__1__18_chany_bottom_out;
wire [0:228] cby_0__1__18_chany_top_out;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__19_ccff_tail;
wire [0:228] cby_0__1__19_chany_bottom_out;
wire [0:228] cby_0__1__19_chany_top_out;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:228] cby_0__1__1_chany_bottom_out;
wire [0:228] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__20_ccff_tail;
wire [0:228] cby_0__1__20_chany_bottom_out;
wire [0:228] cby_0__1__20_chany_top_out;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:228] cby_0__1__2_chany_bottom_out;
wire [0:228] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:228] cby_0__1__3_chany_bottom_out;
wire [0:228] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:228] cby_0__1__4_chany_bottom_out;
wire [0:228] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__5_ccff_tail;
wire [0:228] cby_0__1__5_chany_bottom_out;
wire [0:228] cby_0__1__5_chany_top_out;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__6_ccff_tail;
wire [0:228] cby_0__1__6_chany_bottom_out;
wire [0:228] cby_0__1__6_chany_top_out;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__7_ccff_tail;
wire [0:228] cby_0__1__7_chany_bottom_out;
wire [0:228] cby_0__1__7_chany_top_out;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__8_ccff_tail;
wire [0:228] cby_0__1__8_chany_bottom_out;
wire [0:228] cby_0__1__8_chany_top_out;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__9_ccff_tail;
wire [0:228] cby_0__1__9_chany_bottom_out;
wire [0:228] cby_0__1__9_chany_top_out;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__5__0_ccff_tail;
wire [0:228] cby_0__5__0_chany_bottom_out;
wire [0:228] cby_0__5__0_chany_top_out;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__5__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:228] cby_1__1__0_chany_bottom_out;
wire [0:228] cby_1__1__0_chany_top_out;
wire [0:228] cby_1__1__100_chany_bottom_out;
wire [0:228] cby_1__1__100_chany_top_out;
wire [0:228] cby_1__1__101_chany_bottom_out;
wire [0:228] cby_1__1__101_chany_top_out;
wire [0:228] cby_1__1__102_chany_bottom_out;
wire [0:228] cby_1__1__102_chany_top_out;
wire [0:228] cby_1__1__103_chany_bottom_out;
wire [0:228] cby_1__1__103_chany_top_out;
wire [0:228] cby_1__1__104_chany_bottom_out;
wire [0:228] cby_1__1__104_chany_top_out;
wire [0:228] cby_1__1__105_chany_bottom_out;
wire [0:228] cby_1__1__105_chany_top_out;
wire [0:228] cby_1__1__106_chany_bottom_out;
wire [0:228] cby_1__1__106_chany_top_out;
wire [0:228] cby_1__1__107_chany_bottom_out;
wire [0:228] cby_1__1__107_chany_top_out;
wire [0:228] cby_1__1__108_chany_bottom_out;
wire [0:228] cby_1__1__108_chany_top_out;
wire [0:228] cby_1__1__109_chany_bottom_out;
wire [0:228] cby_1__1__109_chany_top_out;
wire [0:228] cby_1__1__10_chany_bottom_out;
wire [0:228] cby_1__1__10_chany_top_out;
wire [0:228] cby_1__1__110_chany_bottom_out;
wire [0:228] cby_1__1__110_chany_top_out;
wire [0:228] cby_1__1__111_chany_bottom_out;
wire [0:228] cby_1__1__111_chany_top_out;
wire [0:228] cby_1__1__112_chany_bottom_out;
wire [0:228] cby_1__1__112_chany_top_out;
wire [0:228] cby_1__1__113_chany_bottom_out;
wire [0:228] cby_1__1__113_chany_top_out;
wire [0:228] cby_1__1__114_chany_bottom_out;
wire [0:228] cby_1__1__114_chany_top_out;
wire [0:228] cby_1__1__115_chany_bottom_out;
wire [0:228] cby_1__1__115_chany_top_out;
wire [0:228] cby_1__1__116_chany_bottom_out;
wire [0:228] cby_1__1__116_chany_top_out;
wire [0:228] cby_1__1__117_chany_bottom_out;
wire [0:228] cby_1__1__117_chany_top_out;
wire [0:228] cby_1__1__118_chany_bottom_out;
wire [0:228] cby_1__1__118_chany_top_out;
wire [0:228] cby_1__1__119_chany_bottom_out;
wire [0:228] cby_1__1__119_chany_top_out;
wire [0:228] cby_1__1__11_chany_bottom_out;
wire [0:228] cby_1__1__11_chany_top_out;
wire [0:228] cby_1__1__120_chany_bottom_out;
wire [0:228] cby_1__1__120_chany_top_out;
wire [0:228] cby_1__1__121_chany_bottom_out;
wire [0:228] cby_1__1__121_chany_top_out;
wire [0:228] cby_1__1__122_chany_bottom_out;
wire [0:228] cby_1__1__122_chany_top_out;
wire [0:228] cby_1__1__123_chany_bottom_out;
wire [0:228] cby_1__1__123_chany_top_out;
wire [0:228] cby_1__1__124_chany_bottom_out;
wire [0:228] cby_1__1__124_chany_top_out;
wire [0:228] cby_1__1__125_chany_bottom_out;
wire [0:228] cby_1__1__125_chany_top_out;
wire [0:228] cby_1__1__126_chany_bottom_out;
wire [0:228] cby_1__1__126_chany_top_out;
wire [0:228] cby_1__1__127_chany_bottom_out;
wire [0:228] cby_1__1__127_chany_top_out;
wire [0:228] cby_1__1__128_chany_bottom_out;
wire [0:228] cby_1__1__128_chany_top_out;
wire [0:228] cby_1__1__129_chany_bottom_out;
wire [0:228] cby_1__1__129_chany_top_out;
wire [0:228] cby_1__1__12_chany_bottom_out;
wire [0:228] cby_1__1__12_chany_top_out;
wire [0:228] cby_1__1__130_chany_bottom_out;
wire [0:228] cby_1__1__130_chany_top_out;
wire [0:228] cby_1__1__131_chany_bottom_out;
wire [0:228] cby_1__1__131_chany_top_out;
wire [0:228] cby_1__1__132_chany_bottom_out;
wire [0:228] cby_1__1__132_chany_top_out;
wire [0:228] cby_1__1__133_chany_bottom_out;
wire [0:228] cby_1__1__133_chany_top_out;
wire [0:228] cby_1__1__134_chany_bottom_out;
wire [0:228] cby_1__1__134_chany_top_out;
wire [0:228] cby_1__1__135_chany_bottom_out;
wire [0:228] cby_1__1__135_chany_top_out;
wire [0:228] cby_1__1__136_chany_bottom_out;
wire [0:228] cby_1__1__136_chany_top_out;
wire [0:228] cby_1__1__137_chany_bottom_out;
wire [0:228] cby_1__1__137_chany_top_out;
wire [0:228] cby_1__1__138_chany_bottom_out;
wire [0:228] cby_1__1__138_chany_top_out;
wire [0:228] cby_1__1__139_chany_bottom_out;
wire [0:228] cby_1__1__139_chany_top_out;
wire [0:228] cby_1__1__13_chany_bottom_out;
wire [0:228] cby_1__1__13_chany_top_out;
wire [0:228] cby_1__1__140_chany_bottom_out;
wire [0:228] cby_1__1__140_chany_top_out;
wire [0:228] cby_1__1__141_chany_bottom_out;
wire [0:228] cby_1__1__141_chany_top_out;
wire [0:228] cby_1__1__142_chany_bottom_out;
wire [0:228] cby_1__1__142_chany_top_out;
wire [0:228] cby_1__1__143_chany_bottom_out;
wire [0:228] cby_1__1__143_chany_top_out;
wire [0:228] cby_1__1__144_chany_bottom_out;
wire [0:228] cby_1__1__144_chany_top_out;
wire [0:228] cby_1__1__145_chany_bottom_out;
wire [0:228] cby_1__1__145_chany_top_out;
wire [0:228] cby_1__1__146_chany_bottom_out;
wire [0:228] cby_1__1__146_chany_top_out;
wire [0:228] cby_1__1__147_chany_bottom_out;
wire [0:228] cby_1__1__147_chany_top_out;
wire [0:228] cby_1__1__148_chany_bottom_out;
wire [0:228] cby_1__1__148_chany_top_out;
wire [0:228] cby_1__1__149_chany_bottom_out;
wire [0:228] cby_1__1__149_chany_top_out;
wire [0:228] cby_1__1__14_chany_bottom_out;
wire [0:228] cby_1__1__14_chany_top_out;
wire [0:228] cby_1__1__150_chany_bottom_out;
wire [0:228] cby_1__1__150_chany_top_out;
wire [0:228] cby_1__1__151_chany_bottom_out;
wire [0:228] cby_1__1__151_chany_top_out;
wire [0:228] cby_1__1__152_chany_bottom_out;
wire [0:228] cby_1__1__152_chany_top_out;
wire [0:228] cby_1__1__153_chany_bottom_out;
wire [0:228] cby_1__1__153_chany_top_out;
wire [0:228] cby_1__1__154_chany_bottom_out;
wire [0:228] cby_1__1__154_chany_top_out;
wire [0:228] cby_1__1__155_chany_bottom_out;
wire [0:228] cby_1__1__155_chany_top_out;
wire [0:228] cby_1__1__156_chany_bottom_out;
wire [0:228] cby_1__1__156_chany_top_out;
wire [0:228] cby_1__1__157_chany_bottom_out;
wire [0:228] cby_1__1__157_chany_top_out;
wire [0:228] cby_1__1__158_chany_bottom_out;
wire [0:228] cby_1__1__158_chany_top_out;
wire [0:228] cby_1__1__159_chany_bottom_out;
wire [0:228] cby_1__1__159_chany_top_out;
wire [0:228] cby_1__1__15_chany_bottom_out;
wire [0:228] cby_1__1__15_chany_top_out;
wire [0:228] cby_1__1__160_chany_bottom_out;
wire [0:228] cby_1__1__160_chany_top_out;
wire [0:228] cby_1__1__161_chany_bottom_out;
wire [0:228] cby_1__1__161_chany_top_out;
wire [0:228] cby_1__1__162_chany_bottom_out;
wire [0:228] cby_1__1__162_chany_top_out;
wire [0:228] cby_1__1__163_chany_bottom_out;
wire [0:228] cby_1__1__163_chany_top_out;
wire [0:228] cby_1__1__164_chany_bottom_out;
wire [0:228] cby_1__1__164_chany_top_out;
wire [0:228] cby_1__1__165_chany_bottom_out;
wire [0:228] cby_1__1__165_chany_top_out;
wire [0:228] cby_1__1__166_chany_bottom_out;
wire [0:228] cby_1__1__166_chany_top_out;
wire [0:228] cby_1__1__167_chany_bottom_out;
wire [0:228] cby_1__1__167_chany_top_out;
wire [0:228] cby_1__1__168_chany_bottom_out;
wire [0:228] cby_1__1__168_chany_top_out;
wire [0:228] cby_1__1__169_chany_bottom_out;
wire [0:228] cby_1__1__169_chany_top_out;
wire [0:228] cby_1__1__16_chany_bottom_out;
wire [0:228] cby_1__1__16_chany_top_out;
wire [0:228] cby_1__1__170_chany_bottom_out;
wire [0:228] cby_1__1__170_chany_top_out;
wire [0:228] cby_1__1__171_chany_bottom_out;
wire [0:228] cby_1__1__171_chany_top_out;
wire [0:228] cby_1__1__172_chany_bottom_out;
wire [0:228] cby_1__1__172_chany_top_out;
wire [0:228] cby_1__1__173_chany_bottom_out;
wire [0:228] cby_1__1__173_chany_top_out;
wire [0:228] cby_1__1__174_chany_bottom_out;
wire [0:228] cby_1__1__174_chany_top_out;
wire [0:228] cby_1__1__175_chany_bottom_out;
wire [0:228] cby_1__1__175_chany_top_out;
wire [0:228] cby_1__1__176_chany_bottom_out;
wire [0:228] cby_1__1__176_chany_top_out;
wire [0:228] cby_1__1__177_chany_bottom_out;
wire [0:228] cby_1__1__177_chany_top_out;
wire [0:228] cby_1__1__178_chany_bottom_out;
wire [0:228] cby_1__1__178_chany_top_out;
wire [0:228] cby_1__1__179_chany_bottom_out;
wire [0:228] cby_1__1__179_chany_top_out;
wire [0:228] cby_1__1__17_chany_bottom_out;
wire [0:228] cby_1__1__17_chany_top_out;
wire [0:228] cby_1__1__180_chany_bottom_out;
wire [0:228] cby_1__1__180_chany_top_out;
wire [0:228] cby_1__1__181_chany_bottom_out;
wire [0:228] cby_1__1__181_chany_top_out;
wire [0:228] cby_1__1__182_chany_bottom_out;
wire [0:228] cby_1__1__182_chany_top_out;
wire [0:228] cby_1__1__183_chany_bottom_out;
wire [0:228] cby_1__1__183_chany_top_out;
wire [0:228] cby_1__1__184_chany_bottom_out;
wire [0:228] cby_1__1__184_chany_top_out;
wire [0:228] cby_1__1__185_chany_bottom_out;
wire [0:228] cby_1__1__185_chany_top_out;
wire [0:228] cby_1__1__186_chany_bottom_out;
wire [0:228] cby_1__1__186_chany_top_out;
wire [0:228] cby_1__1__187_chany_bottom_out;
wire [0:228] cby_1__1__187_chany_top_out;
wire [0:228] cby_1__1__188_chany_bottom_out;
wire [0:228] cby_1__1__188_chany_top_out;
wire [0:228] cby_1__1__189_chany_bottom_out;
wire [0:228] cby_1__1__189_chany_top_out;
wire [0:228] cby_1__1__18_chany_bottom_out;
wire [0:228] cby_1__1__18_chany_top_out;
wire [0:228] cby_1__1__190_chany_bottom_out;
wire [0:228] cby_1__1__190_chany_top_out;
wire [0:228] cby_1__1__191_chany_bottom_out;
wire [0:228] cby_1__1__191_chany_top_out;
wire [0:228] cby_1__1__192_chany_bottom_out;
wire [0:228] cby_1__1__192_chany_top_out;
wire [0:228] cby_1__1__193_chany_bottom_out;
wire [0:228] cby_1__1__193_chany_top_out;
wire [0:228] cby_1__1__194_chany_bottom_out;
wire [0:228] cby_1__1__194_chany_top_out;
wire [0:228] cby_1__1__195_chany_bottom_out;
wire [0:228] cby_1__1__195_chany_top_out;
wire [0:228] cby_1__1__196_chany_bottom_out;
wire [0:228] cby_1__1__196_chany_top_out;
wire [0:228] cby_1__1__197_chany_bottom_out;
wire [0:228] cby_1__1__197_chany_top_out;
wire [0:228] cby_1__1__198_chany_bottom_out;
wire [0:228] cby_1__1__198_chany_top_out;
wire [0:228] cby_1__1__199_chany_bottom_out;
wire [0:228] cby_1__1__199_chany_top_out;
wire [0:228] cby_1__1__19_chany_bottom_out;
wire [0:228] cby_1__1__19_chany_top_out;
wire [0:228] cby_1__1__1_chany_bottom_out;
wire [0:228] cby_1__1__1_chany_top_out;
wire [0:228] cby_1__1__200_chany_bottom_out;
wire [0:228] cby_1__1__200_chany_top_out;
wire [0:228] cby_1__1__201_chany_bottom_out;
wire [0:228] cby_1__1__201_chany_top_out;
wire [0:228] cby_1__1__202_chany_bottom_out;
wire [0:228] cby_1__1__202_chany_top_out;
wire [0:228] cby_1__1__203_chany_bottom_out;
wire [0:228] cby_1__1__203_chany_top_out;
wire [0:228] cby_1__1__204_chany_bottom_out;
wire [0:228] cby_1__1__204_chany_top_out;
wire [0:228] cby_1__1__205_chany_bottom_out;
wire [0:228] cby_1__1__205_chany_top_out;
wire [0:228] cby_1__1__206_chany_bottom_out;
wire [0:228] cby_1__1__206_chany_top_out;
wire [0:228] cby_1__1__207_chany_bottom_out;
wire [0:228] cby_1__1__207_chany_top_out;
wire [0:228] cby_1__1__208_chany_bottom_out;
wire [0:228] cby_1__1__208_chany_top_out;
wire [0:228] cby_1__1__209_chany_bottom_out;
wire [0:228] cby_1__1__209_chany_top_out;
wire [0:228] cby_1__1__20_chany_bottom_out;
wire [0:228] cby_1__1__20_chany_top_out;
wire [0:228] cby_1__1__210_chany_bottom_out;
wire [0:228] cby_1__1__210_chany_top_out;
wire [0:228] cby_1__1__211_chany_bottom_out;
wire [0:228] cby_1__1__211_chany_top_out;
wire [0:228] cby_1__1__212_chany_bottom_out;
wire [0:228] cby_1__1__212_chany_top_out;
wire [0:228] cby_1__1__213_chany_bottom_out;
wire [0:228] cby_1__1__213_chany_top_out;
wire [0:228] cby_1__1__214_chany_bottom_out;
wire [0:228] cby_1__1__214_chany_top_out;
wire [0:228] cby_1__1__215_chany_bottom_out;
wire [0:228] cby_1__1__215_chany_top_out;
wire [0:228] cby_1__1__216_chany_bottom_out;
wire [0:228] cby_1__1__216_chany_top_out;
wire [0:228] cby_1__1__217_chany_bottom_out;
wire [0:228] cby_1__1__217_chany_top_out;
wire [0:228] cby_1__1__218_chany_bottom_out;
wire [0:228] cby_1__1__218_chany_top_out;
wire [0:228] cby_1__1__219_chany_bottom_out;
wire [0:228] cby_1__1__219_chany_top_out;
wire [0:228] cby_1__1__21_chany_bottom_out;
wire [0:228] cby_1__1__21_chany_top_out;
wire [0:228] cby_1__1__220_chany_bottom_out;
wire [0:228] cby_1__1__220_chany_top_out;
wire [0:228] cby_1__1__221_chany_bottom_out;
wire [0:228] cby_1__1__221_chany_top_out;
wire [0:228] cby_1__1__222_chany_bottom_out;
wire [0:228] cby_1__1__222_chany_top_out;
wire [0:228] cby_1__1__223_chany_bottom_out;
wire [0:228] cby_1__1__223_chany_top_out;
wire [0:228] cby_1__1__224_chany_bottom_out;
wire [0:228] cby_1__1__224_chany_top_out;
wire [0:228] cby_1__1__225_chany_bottom_out;
wire [0:228] cby_1__1__225_chany_top_out;
wire [0:228] cby_1__1__226_chany_bottom_out;
wire [0:228] cby_1__1__226_chany_top_out;
wire [0:228] cby_1__1__227_chany_bottom_out;
wire [0:228] cby_1__1__227_chany_top_out;
wire [0:228] cby_1__1__228_chany_bottom_out;
wire [0:228] cby_1__1__228_chany_top_out;
wire [0:228] cby_1__1__229_chany_bottom_out;
wire [0:228] cby_1__1__229_chany_top_out;
wire [0:228] cby_1__1__22_chany_bottom_out;
wire [0:228] cby_1__1__22_chany_top_out;
wire [0:228] cby_1__1__230_chany_bottom_out;
wire [0:228] cby_1__1__230_chany_top_out;
wire [0:228] cby_1__1__231_chany_bottom_out;
wire [0:228] cby_1__1__231_chany_top_out;
wire [0:228] cby_1__1__232_chany_bottom_out;
wire [0:228] cby_1__1__232_chany_top_out;
wire [0:228] cby_1__1__233_chany_bottom_out;
wire [0:228] cby_1__1__233_chany_top_out;
wire [0:228] cby_1__1__234_chany_bottom_out;
wire [0:228] cby_1__1__234_chany_top_out;
wire [0:228] cby_1__1__235_chany_bottom_out;
wire [0:228] cby_1__1__235_chany_top_out;
wire [0:228] cby_1__1__236_chany_bottom_out;
wire [0:228] cby_1__1__236_chany_top_out;
wire [0:228] cby_1__1__237_chany_bottom_out;
wire [0:228] cby_1__1__237_chany_top_out;
wire [0:228] cby_1__1__238_chany_bottom_out;
wire [0:228] cby_1__1__238_chany_top_out;
wire [0:228] cby_1__1__239_chany_bottom_out;
wire [0:228] cby_1__1__239_chany_top_out;
wire [0:228] cby_1__1__23_chany_bottom_out;
wire [0:228] cby_1__1__23_chany_top_out;
wire [0:228] cby_1__1__240_chany_bottom_out;
wire [0:228] cby_1__1__240_chany_top_out;
wire [0:228] cby_1__1__241_chany_bottom_out;
wire [0:228] cby_1__1__241_chany_top_out;
wire [0:228] cby_1__1__242_chany_bottom_out;
wire [0:228] cby_1__1__242_chany_top_out;
wire [0:228] cby_1__1__243_chany_bottom_out;
wire [0:228] cby_1__1__243_chany_top_out;
wire [0:228] cby_1__1__244_chany_bottom_out;
wire [0:228] cby_1__1__244_chany_top_out;
wire [0:228] cby_1__1__245_chany_bottom_out;
wire [0:228] cby_1__1__245_chany_top_out;
wire [0:228] cby_1__1__246_chany_bottom_out;
wire [0:228] cby_1__1__246_chany_top_out;
wire [0:228] cby_1__1__247_chany_bottom_out;
wire [0:228] cby_1__1__247_chany_top_out;
wire [0:228] cby_1__1__248_chany_bottom_out;
wire [0:228] cby_1__1__248_chany_top_out;
wire [0:228] cby_1__1__249_chany_bottom_out;
wire [0:228] cby_1__1__249_chany_top_out;
wire [0:228] cby_1__1__24_chany_bottom_out;
wire [0:228] cby_1__1__24_chany_top_out;
wire [0:228] cby_1__1__250_chany_bottom_out;
wire [0:228] cby_1__1__250_chany_top_out;
wire [0:228] cby_1__1__251_chany_bottom_out;
wire [0:228] cby_1__1__251_chany_top_out;
wire [0:228] cby_1__1__252_chany_bottom_out;
wire [0:228] cby_1__1__252_chany_top_out;
wire [0:228] cby_1__1__253_chany_bottom_out;
wire [0:228] cby_1__1__253_chany_top_out;
wire [0:228] cby_1__1__254_chany_bottom_out;
wire [0:228] cby_1__1__254_chany_top_out;
wire [0:228] cby_1__1__255_chany_bottom_out;
wire [0:228] cby_1__1__255_chany_top_out;
wire [0:228] cby_1__1__256_chany_bottom_out;
wire [0:228] cby_1__1__256_chany_top_out;
wire [0:228] cby_1__1__257_chany_bottom_out;
wire [0:228] cby_1__1__257_chany_top_out;
wire [0:228] cby_1__1__258_chany_bottom_out;
wire [0:228] cby_1__1__258_chany_top_out;
wire [0:228] cby_1__1__259_chany_bottom_out;
wire [0:228] cby_1__1__259_chany_top_out;
wire [0:228] cby_1__1__25_chany_bottom_out;
wire [0:228] cby_1__1__25_chany_top_out;
wire [0:228] cby_1__1__260_chany_bottom_out;
wire [0:228] cby_1__1__260_chany_top_out;
wire [0:228] cby_1__1__261_chany_bottom_out;
wire [0:228] cby_1__1__261_chany_top_out;
wire [0:228] cby_1__1__262_chany_bottom_out;
wire [0:228] cby_1__1__262_chany_top_out;
wire [0:228] cby_1__1__263_chany_bottom_out;
wire [0:228] cby_1__1__263_chany_top_out;
wire [0:228] cby_1__1__264_chany_bottom_out;
wire [0:228] cby_1__1__264_chany_top_out;
wire [0:228] cby_1__1__265_chany_bottom_out;
wire [0:228] cby_1__1__265_chany_top_out;
wire [0:228] cby_1__1__266_chany_bottom_out;
wire [0:228] cby_1__1__266_chany_top_out;
wire [0:228] cby_1__1__267_chany_bottom_out;
wire [0:228] cby_1__1__267_chany_top_out;
wire [0:228] cby_1__1__268_chany_bottom_out;
wire [0:228] cby_1__1__268_chany_top_out;
wire [0:228] cby_1__1__269_chany_bottom_out;
wire [0:228] cby_1__1__269_chany_top_out;
wire [0:228] cby_1__1__26_chany_bottom_out;
wire [0:228] cby_1__1__26_chany_top_out;
wire [0:228] cby_1__1__270_chany_bottom_out;
wire [0:228] cby_1__1__270_chany_top_out;
wire [0:228] cby_1__1__271_chany_bottom_out;
wire [0:228] cby_1__1__271_chany_top_out;
wire [0:228] cby_1__1__272_chany_bottom_out;
wire [0:228] cby_1__1__272_chany_top_out;
wire [0:228] cby_1__1__273_chany_bottom_out;
wire [0:228] cby_1__1__273_chany_top_out;
wire [0:228] cby_1__1__274_chany_bottom_out;
wire [0:228] cby_1__1__274_chany_top_out;
wire [0:228] cby_1__1__275_chany_bottom_out;
wire [0:228] cby_1__1__275_chany_top_out;
wire [0:228] cby_1__1__276_chany_bottom_out;
wire [0:228] cby_1__1__276_chany_top_out;
wire [0:228] cby_1__1__277_chany_bottom_out;
wire [0:228] cby_1__1__277_chany_top_out;
wire [0:228] cby_1__1__278_chany_bottom_out;
wire [0:228] cby_1__1__278_chany_top_out;
wire [0:228] cby_1__1__279_chany_bottom_out;
wire [0:228] cby_1__1__279_chany_top_out;
wire [0:228] cby_1__1__27_chany_bottom_out;
wire [0:228] cby_1__1__27_chany_top_out;
wire [0:228] cby_1__1__280_chany_bottom_out;
wire [0:228] cby_1__1__280_chany_top_out;
wire [0:228] cby_1__1__281_chany_bottom_out;
wire [0:228] cby_1__1__281_chany_top_out;
wire [0:228] cby_1__1__282_chany_bottom_out;
wire [0:228] cby_1__1__282_chany_top_out;
wire [0:228] cby_1__1__283_chany_bottom_out;
wire [0:228] cby_1__1__283_chany_top_out;
wire [0:228] cby_1__1__284_chany_bottom_out;
wire [0:228] cby_1__1__284_chany_top_out;
wire [0:228] cby_1__1__285_chany_bottom_out;
wire [0:228] cby_1__1__285_chany_top_out;
wire [0:228] cby_1__1__286_chany_bottom_out;
wire [0:228] cby_1__1__286_chany_top_out;
wire [0:228] cby_1__1__287_chany_bottom_out;
wire [0:228] cby_1__1__287_chany_top_out;
wire [0:228] cby_1__1__288_chany_bottom_out;
wire [0:228] cby_1__1__288_chany_top_out;
wire [0:228] cby_1__1__289_chany_bottom_out;
wire [0:228] cby_1__1__289_chany_top_out;
wire [0:228] cby_1__1__28_chany_bottom_out;
wire [0:228] cby_1__1__28_chany_top_out;
wire [0:228] cby_1__1__290_chany_bottom_out;
wire [0:228] cby_1__1__290_chany_top_out;
wire [0:228] cby_1__1__291_chany_bottom_out;
wire [0:228] cby_1__1__291_chany_top_out;
wire [0:228] cby_1__1__292_chany_bottom_out;
wire [0:228] cby_1__1__292_chany_top_out;
wire [0:228] cby_1__1__293_chany_bottom_out;
wire [0:228] cby_1__1__293_chany_top_out;
wire [0:228] cby_1__1__294_chany_bottom_out;
wire [0:228] cby_1__1__294_chany_top_out;
wire [0:228] cby_1__1__295_chany_bottom_out;
wire [0:228] cby_1__1__295_chany_top_out;
wire [0:228] cby_1__1__296_chany_bottom_out;
wire [0:228] cby_1__1__296_chany_top_out;
wire [0:228] cby_1__1__297_chany_bottom_out;
wire [0:228] cby_1__1__297_chany_top_out;
wire [0:228] cby_1__1__298_chany_bottom_out;
wire [0:228] cby_1__1__298_chany_top_out;
wire [0:228] cby_1__1__299_chany_bottom_out;
wire [0:228] cby_1__1__299_chany_top_out;
wire [0:228] cby_1__1__29_chany_bottom_out;
wire [0:228] cby_1__1__29_chany_top_out;
wire [0:228] cby_1__1__2_chany_bottom_out;
wire [0:228] cby_1__1__2_chany_top_out;
wire [0:228] cby_1__1__300_chany_bottom_out;
wire [0:228] cby_1__1__300_chany_top_out;
wire [0:228] cby_1__1__301_chany_bottom_out;
wire [0:228] cby_1__1__301_chany_top_out;
wire [0:228] cby_1__1__302_chany_bottom_out;
wire [0:228] cby_1__1__302_chany_top_out;
wire [0:228] cby_1__1__303_chany_bottom_out;
wire [0:228] cby_1__1__303_chany_top_out;
wire [0:228] cby_1__1__304_chany_bottom_out;
wire [0:228] cby_1__1__304_chany_top_out;
wire [0:228] cby_1__1__305_chany_bottom_out;
wire [0:228] cby_1__1__305_chany_top_out;
wire [0:228] cby_1__1__306_chany_bottom_out;
wire [0:228] cby_1__1__306_chany_top_out;
wire [0:228] cby_1__1__307_chany_bottom_out;
wire [0:228] cby_1__1__307_chany_top_out;
wire [0:228] cby_1__1__308_chany_bottom_out;
wire [0:228] cby_1__1__308_chany_top_out;
wire [0:228] cby_1__1__309_chany_bottom_out;
wire [0:228] cby_1__1__309_chany_top_out;
wire [0:228] cby_1__1__30_chany_bottom_out;
wire [0:228] cby_1__1__30_chany_top_out;
wire [0:228] cby_1__1__310_chany_bottom_out;
wire [0:228] cby_1__1__310_chany_top_out;
wire [0:228] cby_1__1__311_chany_bottom_out;
wire [0:228] cby_1__1__311_chany_top_out;
wire [0:228] cby_1__1__312_chany_bottom_out;
wire [0:228] cby_1__1__312_chany_top_out;
wire [0:228] cby_1__1__313_chany_bottom_out;
wire [0:228] cby_1__1__313_chany_top_out;
wire [0:228] cby_1__1__314_chany_bottom_out;
wire [0:228] cby_1__1__314_chany_top_out;
wire [0:228] cby_1__1__315_chany_bottom_out;
wire [0:228] cby_1__1__315_chany_top_out;
wire [0:228] cby_1__1__316_chany_bottom_out;
wire [0:228] cby_1__1__316_chany_top_out;
wire [0:228] cby_1__1__317_chany_bottom_out;
wire [0:228] cby_1__1__317_chany_top_out;
wire [0:228] cby_1__1__318_chany_bottom_out;
wire [0:228] cby_1__1__318_chany_top_out;
wire [0:228] cby_1__1__319_chany_bottom_out;
wire [0:228] cby_1__1__319_chany_top_out;
wire [0:228] cby_1__1__31_chany_bottom_out;
wire [0:228] cby_1__1__31_chany_top_out;
wire [0:228] cby_1__1__320_chany_bottom_out;
wire [0:228] cby_1__1__320_chany_top_out;
wire [0:228] cby_1__1__321_chany_bottom_out;
wire [0:228] cby_1__1__321_chany_top_out;
wire [0:228] cby_1__1__322_chany_bottom_out;
wire [0:228] cby_1__1__322_chany_top_out;
wire [0:228] cby_1__1__323_chany_bottom_out;
wire [0:228] cby_1__1__323_chany_top_out;
wire [0:228] cby_1__1__324_chany_bottom_out;
wire [0:228] cby_1__1__324_chany_top_out;
wire [0:228] cby_1__1__325_chany_bottom_out;
wire [0:228] cby_1__1__325_chany_top_out;
wire [0:228] cby_1__1__326_chany_bottom_out;
wire [0:228] cby_1__1__326_chany_top_out;
wire [0:228] cby_1__1__327_chany_bottom_out;
wire [0:228] cby_1__1__327_chany_top_out;
wire [0:228] cby_1__1__328_chany_bottom_out;
wire [0:228] cby_1__1__328_chany_top_out;
wire [0:228] cby_1__1__329_chany_bottom_out;
wire [0:228] cby_1__1__329_chany_top_out;
wire [0:228] cby_1__1__32_chany_bottom_out;
wire [0:228] cby_1__1__32_chany_top_out;
wire [0:228] cby_1__1__330_chany_bottom_out;
wire [0:228] cby_1__1__330_chany_top_out;
wire [0:228] cby_1__1__331_chany_bottom_out;
wire [0:228] cby_1__1__331_chany_top_out;
wire [0:228] cby_1__1__332_chany_bottom_out;
wire [0:228] cby_1__1__332_chany_top_out;
wire [0:228] cby_1__1__333_chany_bottom_out;
wire [0:228] cby_1__1__333_chany_top_out;
wire [0:228] cby_1__1__334_chany_bottom_out;
wire [0:228] cby_1__1__334_chany_top_out;
wire [0:228] cby_1__1__335_chany_bottom_out;
wire [0:228] cby_1__1__335_chany_top_out;
wire [0:228] cby_1__1__336_chany_bottom_out;
wire [0:228] cby_1__1__336_chany_top_out;
wire [0:228] cby_1__1__337_chany_bottom_out;
wire [0:228] cby_1__1__337_chany_top_out;
wire [0:228] cby_1__1__338_chany_bottom_out;
wire [0:228] cby_1__1__338_chany_top_out;
wire [0:228] cby_1__1__339_chany_bottom_out;
wire [0:228] cby_1__1__339_chany_top_out;
wire [0:228] cby_1__1__33_chany_bottom_out;
wire [0:228] cby_1__1__33_chany_top_out;
wire [0:228] cby_1__1__340_chany_bottom_out;
wire [0:228] cby_1__1__340_chany_top_out;
wire [0:228] cby_1__1__341_chany_bottom_out;
wire [0:228] cby_1__1__341_chany_top_out;
wire [0:228] cby_1__1__342_chany_bottom_out;
wire [0:228] cby_1__1__342_chany_top_out;
wire [0:228] cby_1__1__343_chany_bottom_out;
wire [0:228] cby_1__1__343_chany_top_out;
wire [0:228] cby_1__1__344_chany_bottom_out;
wire [0:228] cby_1__1__344_chany_top_out;
wire [0:228] cby_1__1__345_chany_bottom_out;
wire [0:228] cby_1__1__345_chany_top_out;
wire [0:228] cby_1__1__346_chany_bottom_out;
wire [0:228] cby_1__1__346_chany_top_out;
wire [0:228] cby_1__1__347_chany_bottom_out;
wire [0:228] cby_1__1__347_chany_top_out;
wire [0:228] cby_1__1__348_chany_bottom_out;
wire [0:228] cby_1__1__348_chany_top_out;
wire [0:228] cby_1__1__349_chany_bottom_out;
wire [0:228] cby_1__1__349_chany_top_out;
wire [0:228] cby_1__1__34_chany_bottom_out;
wire [0:228] cby_1__1__34_chany_top_out;
wire [0:228] cby_1__1__350_chany_bottom_out;
wire [0:228] cby_1__1__350_chany_top_out;
wire [0:228] cby_1__1__351_chany_bottom_out;
wire [0:228] cby_1__1__351_chany_top_out;
wire [0:228] cby_1__1__352_chany_bottom_out;
wire [0:228] cby_1__1__352_chany_top_out;
wire [0:228] cby_1__1__353_chany_bottom_out;
wire [0:228] cby_1__1__353_chany_top_out;
wire [0:228] cby_1__1__354_chany_bottom_out;
wire [0:228] cby_1__1__354_chany_top_out;
wire [0:228] cby_1__1__355_chany_bottom_out;
wire [0:228] cby_1__1__355_chany_top_out;
wire [0:228] cby_1__1__356_chany_bottom_out;
wire [0:228] cby_1__1__356_chany_top_out;
wire [0:228] cby_1__1__357_chany_bottom_out;
wire [0:228] cby_1__1__357_chany_top_out;
wire [0:228] cby_1__1__358_chany_bottom_out;
wire [0:228] cby_1__1__358_chany_top_out;
wire [0:228] cby_1__1__359_chany_bottom_out;
wire [0:228] cby_1__1__359_chany_top_out;
wire [0:228] cby_1__1__35_chany_bottom_out;
wire [0:228] cby_1__1__35_chany_top_out;
wire [0:228] cby_1__1__360_chany_bottom_out;
wire [0:228] cby_1__1__360_chany_top_out;
wire [0:228] cby_1__1__361_chany_bottom_out;
wire [0:228] cby_1__1__361_chany_top_out;
wire [0:228] cby_1__1__362_chany_bottom_out;
wire [0:228] cby_1__1__362_chany_top_out;
wire [0:228] cby_1__1__363_chany_bottom_out;
wire [0:228] cby_1__1__363_chany_top_out;
wire [0:228] cby_1__1__364_chany_bottom_out;
wire [0:228] cby_1__1__364_chany_top_out;
wire [0:228] cby_1__1__365_chany_bottom_out;
wire [0:228] cby_1__1__365_chany_top_out;
wire [0:228] cby_1__1__366_chany_bottom_out;
wire [0:228] cby_1__1__366_chany_top_out;
wire [0:228] cby_1__1__367_chany_bottom_out;
wire [0:228] cby_1__1__367_chany_top_out;
wire [0:228] cby_1__1__368_chany_bottom_out;
wire [0:228] cby_1__1__368_chany_top_out;
wire [0:228] cby_1__1__369_chany_bottom_out;
wire [0:228] cby_1__1__369_chany_top_out;
wire [0:228] cby_1__1__36_chany_bottom_out;
wire [0:228] cby_1__1__36_chany_top_out;
wire [0:228] cby_1__1__370_chany_bottom_out;
wire [0:228] cby_1__1__370_chany_top_out;
wire [0:228] cby_1__1__371_chany_bottom_out;
wire [0:228] cby_1__1__371_chany_top_out;
wire [0:228] cby_1__1__372_chany_bottom_out;
wire [0:228] cby_1__1__372_chany_top_out;
wire [0:228] cby_1__1__373_chany_bottom_out;
wire [0:228] cby_1__1__373_chany_top_out;
wire [0:228] cby_1__1__374_chany_bottom_out;
wire [0:228] cby_1__1__374_chany_top_out;
wire [0:228] cby_1__1__375_chany_bottom_out;
wire [0:228] cby_1__1__375_chany_top_out;
wire [0:228] cby_1__1__376_chany_bottom_out;
wire [0:228] cby_1__1__376_chany_top_out;
wire [0:228] cby_1__1__377_chany_bottom_out;
wire [0:228] cby_1__1__377_chany_top_out;
wire [0:228] cby_1__1__378_chany_bottom_out;
wire [0:228] cby_1__1__378_chany_top_out;
wire [0:228] cby_1__1__379_chany_bottom_out;
wire [0:228] cby_1__1__379_chany_top_out;
wire [0:228] cby_1__1__37_chany_bottom_out;
wire [0:228] cby_1__1__37_chany_top_out;
wire [0:228] cby_1__1__380_chany_bottom_out;
wire [0:228] cby_1__1__380_chany_top_out;
wire [0:228] cby_1__1__381_chany_bottom_out;
wire [0:228] cby_1__1__381_chany_top_out;
wire [0:228] cby_1__1__382_chany_bottom_out;
wire [0:228] cby_1__1__382_chany_top_out;
wire [0:228] cby_1__1__383_chany_bottom_out;
wire [0:228] cby_1__1__383_chany_top_out;
wire [0:228] cby_1__1__384_chany_bottom_out;
wire [0:228] cby_1__1__384_chany_top_out;
wire [0:228] cby_1__1__385_chany_bottom_out;
wire [0:228] cby_1__1__385_chany_top_out;
wire [0:228] cby_1__1__386_chany_bottom_out;
wire [0:228] cby_1__1__386_chany_top_out;
wire [0:228] cby_1__1__387_chany_bottom_out;
wire [0:228] cby_1__1__387_chany_top_out;
wire [0:228] cby_1__1__388_chany_bottom_out;
wire [0:228] cby_1__1__388_chany_top_out;
wire [0:228] cby_1__1__389_chany_bottom_out;
wire [0:228] cby_1__1__389_chany_top_out;
wire [0:228] cby_1__1__38_chany_bottom_out;
wire [0:228] cby_1__1__38_chany_top_out;
wire [0:228] cby_1__1__390_chany_bottom_out;
wire [0:228] cby_1__1__390_chany_top_out;
wire [0:228] cby_1__1__391_chany_bottom_out;
wire [0:228] cby_1__1__391_chany_top_out;
wire [0:228] cby_1__1__392_chany_bottom_out;
wire [0:228] cby_1__1__392_chany_top_out;
wire [0:228] cby_1__1__393_chany_bottom_out;
wire [0:228] cby_1__1__393_chany_top_out;
wire [0:228] cby_1__1__394_chany_bottom_out;
wire [0:228] cby_1__1__394_chany_top_out;
wire [0:228] cby_1__1__395_chany_bottom_out;
wire [0:228] cby_1__1__395_chany_top_out;
wire [0:228] cby_1__1__396_chany_bottom_out;
wire [0:228] cby_1__1__396_chany_top_out;
wire [0:228] cby_1__1__397_chany_bottom_out;
wire [0:228] cby_1__1__397_chany_top_out;
wire [0:228] cby_1__1__398_chany_bottom_out;
wire [0:228] cby_1__1__398_chany_top_out;
wire [0:228] cby_1__1__399_chany_bottom_out;
wire [0:228] cby_1__1__399_chany_top_out;
wire [0:228] cby_1__1__39_chany_bottom_out;
wire [0:228] cby_1__1__39_chany_top_out;
wire [0:228] cby_1__1__3_chany_bottom_out;
wire [0:228] cby_1__1__3_chany_top_out;
wire [0:228] cby_1__1__400_chany_bottom_out;
wire [0:228] cby_1__1__400_chany_top_out;
wire [0:228] cby_1__1__401_chany_bottom_out;
wire [0:228] cby_1__1__401_chany_top_out;
wire [0:228] cby_1__1__402_chany_bottom_out;
wire [0:228] cby_1__1__402_chany_top_out;
wire [0:228] cby_1__1__403_chany_bottom_out;
wire [0:228] cby_1__1__403_chany_top_out;
wire [0:228] cby_1__1__404_chany_bottom_out;
wire [0:228] cby_1__1__404_chany_top_out;
wire [0:228] cby_1__1__405_chany_bottom_out;
wire [0:228] cby_1__1__405_chany_top_out;
wire [0:228] cby_1__1__406_chany_bottom_out;
wire [0:228] cby_1__1__406_chany_top_out;
wire [0:228] cby_1__1__407_chany_bottom_out;
wire [0:228] cby_1__1__407_chany_top_out;
wire [0:228] cby_1__1__408_chany_bottom_out;
wire [0:228] cby_1__1__408_chany_top_out;
wire [0:228] cby_1__1__409_chany_bottom_out;
wire [0:228] cby_1__1__409_chany_top_out;
wire [0:228] cby_1__1__40_chany_bottom_out;
wire [0:228] cby_1__1__40_chany_top_out;
wire [0:228] cby_1__1__410_chany_bottom_out;
wire [0:228] cby_1__1__410_chany_top_out;
wire [0:228] cby_1__1__411_chany_bottom_out;
wire [0:228] cby_1__1__411_chany_top_out;
wire [0:228] cby_1__1__412_chany_bottom_out;
wire [0:228] cby_1__1__412_chany_top_out;
wire [0:228] cby_1__1__413_chany_bottom_out;
wire [0:228] cby_1__1__413_chany_top_out;
wire [0:228] cby_1__1__414_chany_bottom_out;
wire [0:228] cby_1__1__414_chany_top_out;
wire [0:228] cby_1__1__415_chany_bottom_out;
wire [0:228] cby_1__1__415_chany_top_out;
wire [0:228] cby_1__1__416_chany_bottom_out;
wire [0:228] cby_1__1__416_chany_top_out;
wire [0:228] cby_1__1__417_chany_bottom_out;
wire [0:228] cby_1__1__417_chany_top_out;
wire [0:228] cby_1__1__418_chany_bottom_out;
wire [0:228] cby_1__1__418_chany_top_out;
wire [0:228] cby_1__1__419_chany_bottom_out;
wire [0:228] cby_1__1__419_chany_top_out;
wire [0:228] cby_1__1__41_chany_bottom_out;
wire [0:228] cby_1__1__41_chany_top_out;
wire [0:228] cby_1__1__420_chany_bottom_out;
wire [0:228] cby_1__1__420_chany_top_out;
wire [0:228] cby_1__1__421_chany_bottom_out;
wire [0:228] cby_1__1__421_chany_top_out;
wire [0:228] cby_1__1__422_chany_bottom_out;
wire [0:228] cby_1__1__422_chany_top_out;
wire [0:228] cby_1__1__42_chany_bottom_out;
wire [0:228] cby_1__1__42_chany_top_out;
wire [0:228] cby_1__1__43_chany_bottom_out;
wire [0:228] cby_1__1__43_chany_top_out;
wire [0:228] cby_1__1__44_chany_bottom_out;
wire [0:228] cby_1__1__44_chany_top_out;
wire [0:228] cby_1__1__45_chany_bottom_out;
wire [0:228] cby_1__1__45_chany_top_out;
wire [0:228] cby_1__1__46_chany_bottom_out;
wire [0:228] cby_1__1__46_chany_top_out;
wire [0:228] cby_1__1__47_chany_bottom_out;
wire [0:228] cby_1__1__47_chany_top_out;
wire [0:228] cby_1__1__48_chany_bottom_out;
wire [0:228] cby_1__1__48_chany_top_out;
wire [0:228] cby_1__1__49_chany_bottom_out;
wire [0:228] cby_1__1__49_chany_top_out;
wire [0:228] cby_1__1__4_chany_bottom_out;
wire [0:228] cby_1__1__4_chany_top_out;
wire [0:228] cby_1__1__50_chany_bottom_out;
wire [0:228] cby_1__1__50_chany_top_out;
wire [0:228] cby_1__1__51_chany_bottom_out;
wire [0:228] cby_1__1__51_chany_top_out;
wire [0:228] cby_1__1__52_chany_bottom_out;
wire [0:228] cby_1__1__52_chany_top_out;
wire [0:228] cby_1__1__53_chany_bottom_out;
wire [0:228] cby_1__1__53_chany_top_out;
wire [0:228] cby_1__1__54_chany_bottom_out;
wire [0:228] cby_1__1__54_chany_top_out;
wire [0:228] cby_1__1__55_chany_bottom_out;
wire [0:228] cby_1__1__55_chany_top_out;
wire [0:228] cby_1__1__56_chany_bottom_out;
wire [0:228] cby_1__1__56_chany_top_out;
wire [0:228] cby_1__1__57_chany_bottom_out;
wire [0:228] cby_1__1__57_chany_top_out;
wire [0:228] cby_1__1__58_chany_bottom_out;
wire [0:228] cby_1__1__58_chany_top_out;
wire [0:228] cby_1__1__59_chany_bottom_out;
wire [0:228] cby_1__1__59_chany_top_out;
wire [0:228] cby_1__1__5_chany_bottom_out;
wire [0:228] cby_1__1__5_chany_top_out;
wire [0:228] cby_1__1__60_chany_bottom_out;
wire [0:228] cby_1__1__60_chany_top_out;
wire [0:228] cby_1__1__61_chany_bottom_out;
wire [0:228] cby_1__1__61_chany_top_out;
wire [0:228] cby_1__1__62_chany_bottom_out;
wire [0:228] cby_1__1__62_chany_top_out;
wire [0:228] cby_1__1__63_chany_bottom_out;
wire [0:228] cby_1__1__63_chany_top_out;
wire [0:228] cby_1__1__64_chany_bottom_out;
wire [0:228] cby_1__1__64_chany_top_out;
wire [0:228] cby_1__1__65_chany_bottom_out;
wire [0:228] cby_1__1__65_chany_top_out;
wire [0:228] cby_1__1__66_chany_bottom_out;
wire [0:228] cby_1__1__66_chany_top_out;
wire [0:228] cby_1__1__67_chany_bottom_out;
wire [0:228] cby_1__1__67_chany_top_out;
wire [0:228] cby_1__1__68_chany_bottom_out;
wire [0:228] cby_1__1__68_chany_top_out;
wire [0:228] cby_1__1__69_chany_bottom_out;
wire [0:228] cby_1__1__69_chany_top_out;
wire [0:228] cby_1__1__6_chany_bottom_out;
wire [0:228] cby_1__1__6_chany_top_out;
wire [0:228] cby_1__1__70_chany_bottom_out;
wire [0:228] cby_1__1__70_chany_top_out;
wire [0:228] cby_1__1__71_chany_bottom_out;
wire [0:228] cby_1__1__71_chany_top_out;
wire [0:228] cby_1__1__72_chany_bottom_out;
wire [0:228] cby_1__1__72_chany_top_out;
wire [0:228] cby_1__1__73_chany_bottom_out;
wire [0:228] cby_1__1__73_chany_top_out;
wire [0:228] cby_1__1__74_chany_bottom_out;
wire [0:228] cby_1__1__74_chany_top_out;
wire [0:228] cby_1__1__75_chany_bottom_out;
wire [0:228] cby_1__1__75_chany_top_out;
wire [0:228] cby_1__1__76_chany_bottom_out;
wire [0:228] cby_1__1__76_chany_top_out;
wire [0:228] cby_1__1__77_chany_bottom_out;
wire [0:228] cby_1__1__77_chany_top_out;
wire [0:228] cby_1__1__78_chany_bottom_out;
wire [0:228] cby_1__1__78_chany_top_out;
wire [0:228] cby_1__1__79_chany_bottom_out;
wire [0:228] cby_1__1__79_chany_top_out;
wire [0:228] cby_1__1__7_chany_bottom_out;
wire [0:228] cby_1__1__7_chany_top_out;
wire [0:228] cby_1__1__80_chany_bottom_out;
wire [0:228] cby_1__1__80_chany_top_out;
wire [0:228] cby_1__1__81_chany_bottom_out;
wire [0:228] cby_1__1__81_chany_top_out;
wire [0:228] cby_1__1__82_chany_bottom_out;
wire [0:228] cby_1__1__82_chany_top_out;
wire [0:228] cby_1__1__83_chany_bottom_out;
wire [0:228] cby_1__1__83_chany_top_out;
wire [0:228] cby_1__1__84_chany_bottom_out;
wire [0:228] cby_1__1__84_chany_top_out;
wire [0:228] cby_1__1__85_chany_bottom_out;
wire [0:228] cby_1__1__85_chany_top_out;
wire [0:228] cby_1__1__86_chany_bottom_out;
wire [0:228] cby_1__1__86_chany_top_out;
wire [0:228] cby_1__1__87_chany_bottom_out;
wire [0:228] cby_1__1__87_chany_top_out;
wire [0:228] cby_1__1__88_chany_bottom_out;
wire [0:228] cby_1__1__88_chany_top_out;
wire [0:228] cby_1__1__89_chany_bottom_out;
wire [0:228] cby_1__1__89_chany_top_out;
wire [0:228] cby_1__1__8_chany_bottom_out;
wire [0:228] cby_1__1__8_chany_top_out;
wire [0:228] cby_1__1__90_chany_bottom_out;
wire [0:228] cby_1__1__90_chany_top_out;
wire [0:228] cby_1__1__91_chany_bottom_out;
wire [0:228] cby_1__1__91_chany_top_out;
wire [0:228] cby_1__1__92_chany_bottom_out;
wire [0:228] cby_1__1__92_chany_top_out;
wire [0:228] cby_1__1__93_chany_bottom_out;
wire [0:228] cby_1__1__93_chany_top_out;
wire [0:228] cby_1__1__94_chany_bottom_out;
wire [0:228] cby_1__1__94_chany_top_out;
wire [0:228] cby_1__1__95_chany_bottom_out;
wire [0:228] cby_1__1__95_chany_top_out;
wire [0:228] cby_1__1__96_chany_bottom_out;
wire [0:228] cby_1__1__96_chany_top_out;
wire [0:228] cby_1__1__97_chany_bottom_out;
wire [0:228] cby_1__1__97_chany_top_out;
wire [0:228] cby_1__1__98_chany_bottom_out;
wire [0:228] cby_1__1__98_chany_top_out;
wire [0:228] cby_1__1__99_chany_bottom_out;
wire [0:228] cby_1__1__99_chany_top_out;
wire [0:228] cby_1__1__9_chany_bottom_out;
wire [0:228] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__5__0_ccff_tail;
wire [0:228] cby_1__5__0_chany_bottom_out;
wire [0:228] cby_1__5__0_chany_top_out;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__10_ccff_tail;
wire [0:228] cby_1__5__10_chany_bottom_out;
wire [0:228] cby_1__5__10_chany_top_out;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__11_ccff_tail;
wire [0:228] cby_1__5__11_chany_bottom_out;
wire [0:228] cby_1__5__11_chany_top_out;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__12_ccff_tail;
wire [0:228] cby_1__5__12_chany_bottom_out;
wire [0:228] cby_1__5__12_chany_top_out;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__13_ccff_tail;
wire [0:228] cby_1__5__13_chany_bottom_out;
wire [0:228] cby_1__5__13_chany_top_out;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__14_ccff_tail;
wire [0:228] cby_1__5__14_chany_bottom_out;
wire [0:228] cby_1__5__14_chany_top_out;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__15_ccff_tail;
wire [0:228] cby_1__5__15_chany_bottom_out;
wire [0:228] cby_1__5__15_chany_top_out;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__16_ccff_tail;
wire [0:228] cby_1__5__16_chany_bottom_out;
wire [0:228] cby_1__5__16_chany_top_out;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__17_ccff_tail;
wire [0:228] cby_1__5__17_chany_bottom_out;
wire [0:228] cby_1__5__17_chany_top_out;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__18_ccff_tail;
wire [0:228] cby_1__5__18_chany_bottom_out;
wire [0:228] cby_1__5__18_chany_top_out;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__19_ccff_tail;
wire [0:228] cby_1__5__19_chany_bottom_out;
wire [0:228] cby_1__5__19_chany_top_out;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__1_ccff_tail;
wire [0:228] cby_1__5__1_chany_bottom_out;
wire [0:228] cby_1__5__1_chany_top_out;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__20_ccff_tail;
wire [0:228] cby_1__5__20_chany_bottom_out;
wire [0:228] cby_1__5__20_chany_top_out;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__2_ccff_tail;
wire [0:228] cby_1__5__2_chany_bottom_out;
wire [0:228] cby_1__5__2_chany_top_out;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__3_ccff_tail;
wire [0:228] cby_1__5__3_chany_bottom_out;
wire [0:228] cby_1__5__3_chany_top_out;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__4_ccff_tail;
wire [0:228] cby_1__5__4_chany_bottom_out;
wire [0:228] cby_1__5__4_chany_top_out;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__5_ccff_tail;
wire [0:228] cby_1__5__5_chany_bottom_out;
wire [0:228] cby_1__5__5_chany_top_out;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__6_ccff_tail;
wire [0:228] cby_1__5__6_chany_bottom_out;
wire [0:228] cby_1__5__6_chany_top_out;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__7_ccff_tail;
wire [0:228] cby_1__5__7_chany_bottom_out;
wire [0:228] cby_1__5__7_chany_top_out;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__8_ccff_tail;
wire [0:228] cby_1__5__8_chany_bottom_out;
wire [0:228] cby_1__5__8_chany_top_out;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__5__9_ccff_tail;
wire [0:228] cby_1__5__9_chany_bottom_out;
wire [0:228] cby_1__5__9_chany_top_out;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_22__1__0_ccff_tail;
wire [0:228] cby_22__1__0_chany_bottom_out;
wire [0:228] cby_22__1__0_chany_top_out;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__10_ccff_tail;
wire [0:228] cby_22__1__10_chany_bottom_out;
wire [0:228] cby_22__1__10_chany_top_out;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__11_ccff_tail;
wire [0:228] cby_22__1__11_chany_bottom_out;
wire [0:228] cby_22__1__11_chany_top_out;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__12_ccff_tail;
wire [0:228] cby_22__1__12_chany_bottom_out;
wire [0:228] cby_22__1__12_chany_top_out;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__13_ccff_tail;
wire [0:228] cby_22__1__13_chany_bottom_out;
wire [0:228] cby_22__1__13_chany_top_out;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__14_ccff_tail;
wire [0:228] cby_22__1__14_chany_bottom_out;
wire [0:228] cby_22__1__14_chany_top_out;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__15_ccff_tail;
wire [0:228] cby_22__1__15_chany_bottom_out;
wire [0:228] cby_22__1__15_chany_top_out;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__16_ccff_tail;
wire [0:228] cby_22__1__16_chany_bottom_out;
wire [0:228] cby_22__1__16_chany_top_out;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__17_ccff_tail;
wire [0:228] cby_22__1__17_chany_bottom_out;
wire [0:228] cby_22__1__17_chany_top_out;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__18_ccff_tail;
wire [0:228] cby_22__1__18_chany_bottom_out;
wire [0:228] cby_22__1__18_chany_top_out;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__19_ccff_tail;
wire [0:228] cby_22__1__19_chany_bottom_out;
wire [0:228] cby_22__1__19_chany_top_out;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__1_ccff_tail;
wire [0:228] cby_22__1__1_chany_bottom_out;
wire [0:228] cby_22__1__1_chany_top_out;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__20_ccff_tail;
wire [0:228] cby_22__1__20_chany_bottom_out;
wire [0:228] cby_22__1__20_chany_top_out;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__2_ccff_tail;
wire [0:228] cby_22__1__2_chany_bottom_out;
wire [0:228] cby_22__1__2_chany_top_out;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__3_ccff_tail;
wire [0:228] cby_22__1__3_chany_bottom_out;
wire [0:228] cby_22__1__3_chany_top_out;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__4_ccff_tail;
wire [0:228] cby_22__1__4_chany_bottom_out;
wire [0:228] cby_22__1__4_chany_top_out;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__5_ccff_tail;
wire [0:228] cby_22__1__5_chany_bottom_out;
wire [0:228] cby_22__1__5_chany_top_out;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__6_ccff_tail;
wire [0:228] cby_22__1__6_chany_bottom_out;
wire [0:228] cby_22__1__6_chany_top_out;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__7_ccff_tail;
wire [0:228] cby_22__1__7_chany_bottom_out;
wire [0:228] cby_22__1__7_chany_top_out;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__8_ccff_tail;
wire [0:228] cby_22__1__8_chany_bottom_out;
wire [0:228] cby_22__1__8_chany_top_out;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__1__9_ccff_tail;
wire [0:228] cby_22__1__9_chany_bottom_out;
wire [0:228] cby_22__1__9_chany_top_out;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_22__5__0_ccff_tail;
wire [0:228] cby_22__5__0_chany_bottom_out;
wire [0:228] cby_22__5__0_chany_top_out;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_22__5__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_2__3__0_ccff_tail;
wire [0:228] cby_2__3__0_chany_bottom_out;
wire [0:228] cby_2__3__0_chany_top_out;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__1_ccff_tail;
wire [0:228] cby_2__3__1_chany_bottom_out;
wire [0:228] cby_2__3__1_chany_top_out;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__2_ccff_tail;
wire [0:228] cby_2__3__2_chany_bottom_out;
wire [0:228] cby_2__3__2_chany_top_out;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__3_ccff_tail;
wire [0:228] cby_2__3__3_chany_bottom_out;
wire [0:228] cby_2__3__3_chany_top_out;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__4_ccff_tail;
wire [0:228] cby_2__3__4_chany_bottom_out;
wire [0:228] cby_2__3__4_chany_top_out;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__5_ccff_tail;
wire [0:228] cby_2__3__5_chany_bottom_out;
wire [0:228] cby_2__3__5_chany_top_out;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__6_ccff_tail;
wire [0:228] cby_2__3__6_chany_bottom_out;
wire [0:228] cby_2__3__6_chany_top_out;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__7_ccff_tail;
wire [0:228] cby_2__3__7_chany_bottom_out;
wire [0:228] cby_2__3__7_chany_top_out;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_2__3__8_ccff_tail;
wire [0:228] cby_2__3__8_chany_bottom_out;
wire [0:228] cby_2__3__8_chany_top_out;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cby_3__3__0_ccff_tail;
wire [0:228] cby_3__3__0_chany_bottom_out;
wire [0:228] cby_3__3__0_chany_top_out;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__1_ccff_tail;
wire [0:228] cby_3__3__1_chany_bottom_out;
wire [0:228] cby_3__3__1_chany_top_out;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__2_ccff_tail;
wire [0:228] cby_3__3__2_chany_bottom_out;
wire [0:228] cby_3__3__2_chany_top_out;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__3_ccff_tail;
wire [0:228] cby_3__3__3_chany_bottom_out;
wire [0:228] cby_3__3__3_chany_top_out;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__4_ccff_tail;
wire [0:228] cby_3__3__4_chany_bottom_out;
wire [0:228] cby_3__3__4_chany_top_out;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__5_ccff_tail;
wire [0:228] cby_3__3__5_chany_bottom_out;
wire [0:228] cby_3__3__5_chany_top_out;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__6_ccff_tail;
wire [0:228] cby_3__3__6_chany_bottom_out;
wire [0:228] cby_3__3__6_chany_top_out;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__7_ccff_tail;
wire [0:228] cby_3__3__7_chany_bottom_out;
wire [0:228] cby_3__3__7_chany_top_out;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cby_3__3__8_ccff_tail;
wire [0:228] cby_3__3__8_chany_bottom_out;
wire [0:228] cby_3__3__8_chany_top_out;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_10__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_11__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_12__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_13__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_14__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_15__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_16__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_17__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_18__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_19__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_20__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_21__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_22__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_6__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_7__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_8__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_9__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_ccff_tail;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_ccff_tail;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_ccff_tail;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_ccff_tail;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_ccff_tail;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_14_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_ccff_tail;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_15_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_ccff_tail;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_16_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_ccff_tail;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_17_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_ccff_tail;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_18_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_ccff_tail;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_19_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_ccff_tail;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_20_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_ccff_tail;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_21_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_ccff_tail;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_ccff_tail;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_ccff_tail;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_ccff_tail;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_10_ccff_tail;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_10_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_11_ccff_tail;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_11_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_12_ccff_tail;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_12_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_13_ccff_tail;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_13_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_14_ccff_tail;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_14_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_15_ccff_tail;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_15_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_16_ccff_tail;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_16_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_17_ccff_tail;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_17_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_18_ccff_tail;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_18_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_19_ccff_tail;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_19_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_20_ccff_tail;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_20_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_21_ccff_tail;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_21_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_2_ccff_tail;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_3_ccff_tail;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_4_ccff_tail;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_5_ccff_tail;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_6_ccff_tail;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_7_ccff_tail;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_8_ccff_tail;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_9_ccff_tail;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_10_ccff_tail;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_10_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_11_ccff_tail;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_11_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_12_ccff_tail;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_12_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_13_ccff_tail;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_13_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_14_ccff_tail;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_14_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_15_ccff_tail;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_15_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_16_ccff_tail;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_16_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_17_ccff_tail;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_17_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_18_ccff_tail;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_18_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_19_ccff_tail;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_19_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_20_ccff_tail;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_20_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_21_ccff_tail;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_21_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_2_ccff_tail;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_3_ccff_tail;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_4_ccff_tail;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_5_ccff_tail;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_6_ccff_tail;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_7_ccff_tail;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8_ccff_tail;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_9_ccff_tail;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_10_ccff_tail;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_11_ccff_tail;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_12_ccff_tail;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_13_ccff_tail;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_14_ccff_tail;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_15_ccff_tail;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_16_ccff_tail;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_17_ccff_tail;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_18_ccff_tail;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_19_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_20_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_20_ccff_tail;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_21_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_21_ccff_tail;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_2_ccff_tail;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_3_ccff_tail;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_4_ccff_tail;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_5_ccff_tail;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_6_ccff_tail;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_7_ccff_tail;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_8_ccff_tail;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_9_ccff_tail;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_3__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_3__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_3__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_4_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_4_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_5_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_5_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_6__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_6__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_6_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_6_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_7_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_7_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_8_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_8_top_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_9__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_9__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_9__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:228] sb_0__0__0_chanx_right_out;
wire [0:228] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:228] sb_0__1__0_chanx_right_out;
wire [0:228] sb_0__1__0_chany_bottom_out;
wire [0:228] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__10_ccff_tail;
wire [0:228] sb_0__1__10_chanx_right_out;
wire [0:228] sb_0__1__10_chany_bottom_out;
wire [0:228] sb_0__1__10_chany_top_out;
wire [0:0] sb_0__1__11_ccff_tail;
wire [0:228] sb_0__1__11_chanx_right_out;
wire [0:228] sb_0__1__11_chany_bottom_out;
wire [0:228] sb_0__1__11_chany_top_out;
wire [0:0] sb_0__1__12_ccff_tail;
wire [0:228] sb_0__1__12_chanx_right_out;
wire [0:228] sb_0__1__12_chany_bottom_out;
wire [0:228] sb_0__1__12_chany_top_out;
wire [0:0] sb_0__1__13_ccff_tail;
wire [0:228] sb_0__1__13_chanx_right_out;
wire [0:228] sb_0__1__13_chany_bottom_out;
wire [0:228] sb_0__1__13_chany_top_out;
wire [0:0] sb_0__1__14_ccff_tail;
wire [0:228] sb_0__1__14_chanx_right_out;
wire [0:228] sb_0__1__14_chany_bottom_out;
wire [0:228] sb_0__1__14_chany_top_out;
wire [0:0] sb_0__1__15_ccff_tail;
wire [0:228] sb_0__1__15_chanx_right_out;
wire [0:228] sb_0__1__15_chany_bottom_out;
wire [0:228] sb_0__1__15_chany_top_out;
wire [0:0] sb_0__1__16_ccff_tail;
wire [0:228] sb_0__1__16_chanx_right_out;
wire [0:228] sb_0__1__16_chany_bottom_out;
wire [0:228] sb_0__1__16_chany_top_out;
wire [0:0] sb_0__1__17_ccff_tail;
wire [0:228] sb_0__1__17_chanx_right_out;
wire [0:228] sb_0__1__17_chany_bottom_out;
wire [0:228] sb_0__1__17_chany_top_out;
wire [0:0] sb_0__1__18_ccff_tail;
wire [0:228] sb_0__1__18_chanx_right_out;
wire [0:228] sb_0__1__18_chany_bottom_out;
wire [0:228] sb_0__1__18_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:228] sb_0__1__1_chanx_right_out;
wire [0:228] sb_0__1__1_chany_bottom_out;
wire [0:228] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__1__2_ccff_tail;
wire [0:228] sb_0__1__2_chanx_right_out;
wire [0:228] sb_0__1__2_chany_bottom_out;
wire [0:228] sb_0__1__2_chany_top_out;
wire [0:0] sb_0__1__3_ccff_tail;
wire [0:228] sb_0__1__3_chanx_right_out;
wire [0:228] sb_0__1__3_chany_bottom_out;
wire [0:228] sb_0__1__3_chany_top_out;
wire [0:0] sb_0__1__4_ccff_tail;
wire [0:228] sb_0__1__4_chanx_right_out;
wire [0:228] sb_0__1__4_chany_bottom_out;
wire [0:228] sb_0__1__4_chany_top_out;
wire [0:0] sb_0__1__5_ccff_tail;
wire [0:228] sb_0__1__5_chanx_right_out;
wire [0:228] sb_0__1__5_chany_bottom_out;
wire [0:228] sb_0__1__5_chany_top_out;
wire [0:0] sb_0__1__6_ccff_tail;
wire [0:228] sb_0__1__6_chanx_right_out;
wire [0:228] sb_0__1__6_chany_bottom_out;
wire [0:228] sb_0__1__6_chany_top_out;
wire [0:0] sb_0__1__7_ccff_tail;
wire [0:228] sb_0__1__7_chanx_right_out;
wire [0:228] sb_0__1__7_chany_bottom_out;
wire [0:228] sb_0__1__7_chany_top_out;
wire [0:0] sb_0__1__8_ccff_tail;
wire [0:228] sb_0__1__8_chanx_right_out;
wire [0:228] sb_0__1__8_chany_bottom_out;
wire [0:228] sb_0__1__8_chany_top_out;
wire [0:0] sb_0__1__9_ccff_tail;
wire [0:228] sb_0__1__9_chanx_right_out;
wire [0:228] sb_0__1__9_chany_bottom_out;
wire [0:228] sb_0__1__9_chany_top_out;
wire [0:0] sb_0__22__0_ccff_tail;
wire [0:228] sb_0__22__0_chanx_right_out;
wire [0:228] sb_0__22__0_chany_bottom_out;
wire [0:0] sb_0__4__0_ccff_tail;
wire [0:228] sb_0__4__0_chanx_right_out;
wire [0:228] sb_0__4__0_chany_bottom_out;
wire [0:228] sb_0__4__0_chany_top_out;
wire [0:0] sb_0__5__0_ccff_tail;
wire [0:228] sb_0__5__0_chanx_right_out;
wire [0:228] sb_0__5__0_chany_bottom_out;
wire [0:228] sb_0__5__0_chany_top_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:228] sb_1__0__0_chanx_left_out;
wire [0:228] sb_1__0__0_chanx_right_out;
wire [0:228] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__10_ccff_tail;
wire [0:228] sb_1__0__10_chanx_left_out;
wire [0:228] sb_1__0__10_chanx_right_out;
wire [0:228] sb_1__0__10_chany_top_out;
wire [0:0] sb_1__0__11_ccff_tail;
wire [0:228] sb_1__0__11_chanx_left_out;
wire [0:228] sb_1__0__11_chanx_right_out;
wire [0:228] sb_1__0__11_chany_top_out;
wire [0:0] sb_1__0__12_ccff_tail;
wire [0:228] sb_1__0__12_chanx_left_out;
wire [0:228] sb_1__0__12_chanx_right_out;
wire [0:228] sb_1__0__12_chany_top_out;
wire [0:0] sb_1__0__13_ccff_tail;
wire [0:228] sb_1__0__13_chanx_left_out;
wire [0:228] sb_1__0__13_chanx_right_out;
wire [0:228] sb_1__0__13_chany_top_out;
wire [0:0] sb_1__0__14_ccff_tail;
wire [0:228] sb_1__0__14_chanx_left_out;
wire [0:228] sb_1__0__14_chanx_right_out;
wire [0:228] sb_1__0__14_chany_top_out;
wire [0:0] sb_1__0__15_ccff_tail;
wire [0:228] sb_1__0__15_chanx_left_out;
wire [0:228] sb_1__0__15_chanx_right_out;
wire [0:228] sb_1__0__15_chany_top_out;
wire [0:0] sb_1__0__16_ccff_tail;
wire [0:228] sb_1__0__16_chanx_left_out;
wire [0:228] sb_1__0__16_chanx_right_out;
wire [0:228] sb_1__0__16_chany_top_out;
wire [0:0] sb_1__0__17_ccff_tail;
wire [0:228] sb_1__0__17_chanx_left_out;
wire [0:228] sb_1__0__17_chanx_right_out;
wire [0:228] sb_1__0__17_chany_top_out;
wire [0:0] sb_1__0__18_ccff_tail;
wire [0:228] sb_1__0__18_chanx_left_out;
wire [0:228] sb_1__0__18_chanx_right_out;
wire [0:228] sb_1__0__18_chany_top_out;
wire [0:0] sb_1__0__19_ccff_tail;
wire [0:228] sb_1__0__19_chanx_left_out;
wire [0:228] sb_1__0__19_chanx_right_out;
wire [0:228] sb_1__0__19_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:228] sb_1__0__1_chanx_left_out;
wire [0:228] sb_1__0__1_chanx_right_out;
wire [0:228] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__20_ccff_tail;
wire [0:228] sb_1__0__20_chanx_left_out;
wire [0:228] sb_1__0__20_chanx_right_out;
wire [0:228] sb_1__0__20_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:228] sb_1__0__2_chanx_left_out;
wire [0:228] sb_1__0__2_chanx_right_out;
wire [0:228] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:228] sb_1__0__3_chanx_left_out;
wire [0:228] sb_1__0__3_chanx_right_out;
wire [0:228] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:228] sb_1__0__4_chanx_left_out;
wire [0:228] sb_1__0__4_chanx_right_out;
wire [0:228] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__0__5_ccff_tail;
wire [0:228] sb_1__0__5_chanx_left_out;
wire [0:228] sb_1__0__5_chanx_right_out;
wire [0:228] sb_1__0__5_chany_top_out;
wire [0:0] sb_1__0__6_ccff_tail;
wire [0:228] sb_1__0__6_chanx_left_out;
wire [0:228] sb_1__0__6_chanx_right_out;
wire [0:228] sb_1__0__6_chany_top_out;
wire [0:0] sb_1__0__7_ccff_tail;
wire [0:228] sb_1__0__7_chanx_left_out;
wire [0:228] sb_1__0__7_chanx_right_out;
wire [0:228] sb_1__0__7_chany_top_out;
wire [0:0] sb_1__0__8_ccff_tail;
wire [0:228] sb_1__0__8_chanx_left_out;
wire [0:228] sb_1__0__8_chanx_right_out;
wire [0:228] sb_1__0__8_chany_top_out;
wire [0:0] sb_1__0__9_ccff_tail;
wire [0:228] sb_1__0__9_chanx_left_out;
wire [0:228] sb_1__0__9_chanx_right_out;
wire [0:228] sb_1__0__9_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:228] sb_1__1__0_chanx_left_out;
wire [0:228] sb_1__1__0_chanx_right_out;
wire [0:228] sb_1__1__0_chany_bottom_out;
wire [0:228] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__100_ccff_tail;
wire [0:228] sb_1__1__100_chanx_left_out;
wire [0:228] sb_1__1__100_chanx_right_out;
wire [0:228] sb_1__1__100_chany_bottom_out;
wire [0:228] sb_1__1__100_chany_top_out;
wire [0:0] sb_1__1__101_ccff_tail;
wire [0:228] sb_1__1__101_chanx_left_out;
wire [0:228] sb_1__1__101_chanx_right_out;
wire [0:228] sb_1__1__101_chany_bottom_out;
wire [0:228] sb_1__1__101_chany_top_out;
wire [0:0] sb_1__1__102_ccff_tail;
wire [0:228] sb_1__1__102_chanx_left_out;
wire [0:228] sb_1__1__102_chanx_right_out;
wire [0:228] sb_1__1__102_chany_bottom_out;
wire [0:228] sb_1__1__102_chany_top_out;
wire [0:0] sb_1__1__103_ccff_tail;
wire [0:228] sb_1__1__103_chanx_left_out;
wire [0:228] sb_1__1__103_chanx_right_out;
wire [0:228] sb_1__1__103_chany_bottom_out;
wire [0:228] sb_1__1__103_chany_top_out;
wire [0:0] sb_1__1__104_ccff_tail;
wire [0:228] sb_1__1__104_chanx_left_out;
wire [0:228] sb_1__1__104_chanx_right_out;
wire [0:228] sb_1__1__104_chany_bottom_out;
wire [0:228] sb_1__1__104_chany_top_out;
wire [0:0] sb_1__1__105_ccff_tail;
wire [0:228] sb_1__1__105_chanx_left_out;
wire [0:228] sb_1__1__105_chanx_right_out;
wire [0:228] sb_1__1__105_chany_bottom_out;
wire [0:228] sb_1__1__105_chany_top_out;
wire [0:0] sb_1__1__106_ccff_tail;
wire [0:228] sb_1__1__106_chanx_left_out;
wire [0:228] sb_1__1__106_chanx_right_out;
wire [0:228] sb_1__1__106_chany_bottom_out;
wire [0:228] sb_1__1__106_chany_top_out;
wire [0:0] sb_1__1__107_ccff_tail;
wire [0:228] sb_1__1__107_chanx_left_out;
wire [0:228] sb_1__1__107_chanx_right_out;
wire [0:228] sb_1__1__107_chany_bottom_out;
wire [0:228] sb_1__1__107_chany_top_out;
wire [0:0] sb_1__1__108_ccff_tail;
wire [0:228] sb_1__1__108_chanx_left_out;
wire [0:228] sb_1__1__108_chanx_right_out;
wire [0:228] sb_1__1__108_chany_bottom_out;
wire [0:228] sb_1__1__108_chany_top_out;
wire [0:0] sb_1__1__109_ccff_tail;
wire [0:228] sb_1__1__109_chanx_left_out;
wire [0:228] sb_1__1__109_chanx_right_out;
wire [0:228] sb_1__1__109_chany_bottom_out;
wire [0:228] sb_1__1__109_chany_top_out;
wire [0:0] sb_1__1__10_ccff_tail;
wire [0:228] sb_1__1__10_chanx_left_out;
wire [0:228] sb_1__1__10_chanx_right_out;
wire [0:228] sb_1__1__10_chany_bottom_out;
wire [0:228] sb_1__1__10_chany_top_out;
wire [0:0] sb_1__1__110_ccff_tail;
wire [0:228] sb_1__1__110_chanx_left_out;
wire [0:228] sb_1__1__110_chanx_right_out;
wire [0:228] sb_1__1__110_chany_bottom_out;
wire [0:228] sb_1__1__110_chany_top_out;
wire [0:0] sb_1__1__111_ccff_tail;
wire [0:228] sb_1__1__111_chanx_left_out;
wire [0:228] sb_1__1__111_chanx_right_out;
wire [0:228] sb_1__1__111_chany_bottom_out;
wire [0:228] sb_1__1__111_chany_top_out;
wire [0:0] sb_1__1__112_ccff_tail;
wire [0:228] sb_1__1__112_chanx_left_out;
wire [0:228] sb_1__1__112_chanx_right_out;
wire [0:228] sb_1__1__112_chany_bottom_out;
wire [0:228] sb_1__1__112_chany_top_out;
wire [0:0] sb_1__1__113_ccff_tail;
wire [0:228] sb_1__1__113_chanx_left_out;
wire [0:228] sb_1__1__113_chanx_right_out;
wire [0:228] sb_1__1__113_chany_bottom_out;
wire [0:228] sb_1__1__113_chany_top_out;
wire [0:0] sb_1__1__114_ccff_tail;
wire [0:228] sb_1__1__114_chanx_left_out;
wire [0:228] sb_1__1__114_chanx_right_out;
wire [0:228] sb_1__1__114_chany_bottom_out;
wire [0:228] sb_1__1__114_chany_top_out;
wire [0:0] sb_1__1__115_ccff_tail;
wire [0:228] sb_1__1__115_chanx_left_out;
wire [0:228] sb_1__1__115_chanx_right_out;
wire [0:228] sb_1__1__115_chany_bottom_out;
wire [0:228] sb_1__1__115_chany_top_out;
wire [0:0] sb_1__1__116_ccff_tail;
wire [0:228] sb_1__1__116_chanx_left_out;
wire [0:228] sb_1__1__116_chanx_right_out;
wire [0:228] sb_1__1__116_chany_bottom_out;
wire [0:228] sb_1__1__116_chany_top_out;
wire [0:0] sb_1__1__117_ccff_tail;
wire [0:228] sb_1__1__117_chanx_left_out;
wire [0:228] sb_1__1__117_chanx_right_out;
wire [0:228] sb_1__1__117_chany_bottom_out;
wire [0:228] sb_1__1__117_chany_top_out;
wire [0:0] sb_1__1__118_ccff_tail;
wire [0:228] sb_1__1__118_chanx_left_out;
wire [0:228] sb_1__1__118_chanx_right_out;
wire [0:228] sb_1__1__118_chany_bottom_out;
wire [0:228] sb_1__1__118_chany_top_out;
wire [0:0] sb_1__1__119_ccff_tail;
wire [0:228] sb_1__1__119_chanx_left_out;
wire [0:228] sb_1__1__119_chanx_right_out;
wire [0:228] sb_1__1__119_chany_bottom_out;
wire [0:228] sb_1__1__119_chany_top_out;
wire [0:0] sb_1__1__11_ccff_tail;
wire [0:228] sb_1__1__11_chanx_left_out;
wire [0:228] sb_1__1__11_chanx_right_out;
wire [0:228] sb_1__1__11_chany_bottom_out;
wire [0:228] sb_1__1__11_chany_top_out;
wire [0:0] sb_1__1__120_ccff_tail;
wire [0:228] sb_1__1__120_chanx_left_out;
wire [0:228] sb_1__1__120_chanx_right_out;
wire [0:228] sb_1__1__120_chany_bottom_out;
wire [0:228] sb_1__1__120_chany_top_out;
wire [0:0] sb_1__1__121_ccff_tail;
wire [0:228] sb_1__1__121_chanx_left_out;
wire [0:228] sb_1__1__121_chanx_right_out;
wire [0:228] sb_1__1__121_chany_bottom_out;
wire [0:228] sb_1__1__121_chany_top_out;
wire [0:0] sb_1__1__122_ccff_tail;
wire [0:228] sb_1__1__122_chanx_left_out;
wire [0:228] sb_1__1__122_chanx_right_out;
wire [0:228] sb_1__1__122_chany_bottom_out;
wire [0:228] sb_1__1__122_chany_top_out;
wire [0:0] sb_1__1__123_ccff_tail;
wire [0:228] sb_1__1__123_chanx_left_out;
wire [0:228] sb_1__1__123_chanx_right_out;
wire [0:228] sb_1__1__123_chany_bottom_out;
wire [0:228] sb_1__1__123_chany_top_out;
wire [0:0] sb_1__1__124_ccff_tail;
wire [0:228] sb_1__1__124_chanx_left_out;
wire [0:228] sb_1__1__124_chanx_right_out;
wire [0:228] sb_1__1__124_chany_bottom_out;
wire [0:228] sb_1__1__124_chany_top_out;
wire [0:0] sb_1__1__125_ccff_tail;
wire [0:228] sb_1__1__125_chanx_left_out;
wire [0:228] sb_1__1__125_chanx_right_out;
wire [0:228] sb_1__1__125_chany_bottom_out;
wire [0:228] sb_1__1__125_chany_top_out;
wire [0:0] sb_1__1__126_ccff_tail;
wire [0:228] sb_1__1__126_chanx_left_out;
wire [0:228] sb_1__1__126_chanx_right_out;
wire [0:228] sb_1__1__126_chany_bottom_out;
wire [0:228] sb_1__1__126_chany_top_out;
wire [0:0] sb_1__1__127_ccff_tail;
wire [0:228] sb_1__1__127_chanx_left_out;
wire [0:228] sb_1__1__127_chanx_right_out;
wire [0:228] sb_1__1__127_chany_bottom_out;
wire [0:228] sb_1__1__127_chany_top_out;
wire [0:0] sb_1__1__128_ccff_tail;
wire [0:228] sb_1__1__128_chanx_left_out;
wire [0:228] sb_1__1__128_chanx_right_out;
wire [0:228] sb_1__1__128_chany_bottom_out;
wire [0:228] sb_1__1__128_chany_top_out;
wire [0:0] sb_1__1__129_ccff_tail;
wire [0:228] sb_1__1__129_chanx_left_out;
wire [0:228] sb_1__1__129_chanx_right_out;
wire [0:228] sb_1__1__129_chany_bottom_out;
wire [0:228] sb_1__1__129_chany_top_out;
wire [0:0] sb_1__1__12_ccff_tail;
wire [0:228] sb_1__1__12_chanx_left_out;
wire [0:228] sb_1__1__12_chanx_right_out;
wire [0:228] sb_1__1__12_chany_bottom_out;
wire [0:228] sb_1__1__12_chany_top_out;
wire [0:0] sb_1__1__130_ccff_tail;
wire [0:228] sb_1__1__130_chanx_left_out;
wire [0:228] sb_1__1__130_chanx_right_out;
wire [0:228] sb_1__1__130_chany_bottom_out;
wire [0:228] sb_1__1__130_chany_top_out;
wire [0:0] sb_1__1__131_ccff_tail;
wire [0:228] sb_1__1__131_chanx_left_out;
wire [0:228] sb_1__1__131_chanx_right_out;
wire [0:228] sb_1__1__131_chany_bottom_out;
wire [0:228] sb_1__1__131_chany_top_out;
wire [0:0] sb_1__1__132_ccff_tail;
wire [0:228] sb_1__1__132_chanx_left_out;
wire [0:228] sb_1__1__132_chanx_right_out;
wire [0:228] sb_1__1__132_chany_bottom_out;
wire [0:228] sb_1__1__132_chany_top_out;
wire [0:0] sb_1__1__133_ccff_tail;
wire [0:228] sb_1__1__133_chanx_left_out;
wire [0:228] sb_1__1__133_chanx_right_out;
wire [0:228] sb_1__1__133_chany_bottom_out;
wire [0:228] sb_1__1__133_chany_top_out;
wire [0:0] sb_1__1__134_ccff_tail;
wire [0:228] sb_1__1__134_chanx_left_out;
wire [0:228] sb_1__1__134_chanx_right_out;
wire [0:228] sb_1__1__134_chany_bottom_out;
wire [0:228] sb_1__1__134_chany_top_out;
wire [0:0] sb_1__1__135_ccff_tail;
wire [0:228] sb_1__1__135_chanx_left_out;
wire [0:228] sb_1__1__135_chanx_right_out;
wire [0:228] sb_1__1__135_chany_bottom_out;
wire [0:228] sb_1__1__135_chany_top_out;
wire [0:0] sb_1__1__136_ccff_tail;
wire [0:228] sb_1__1__136_chanx_left_out;
wire [0:228] sb_1__1__136_chanx_right_out;
wire [0:228] sb_1__1__136_chany_bottom_out;
wire [0:228] sb_1__1__136_chany_top_out;
wire [0:0] sb_1__1__137_ccff_tail;
wire [0:228] sb_1__1__137_chanx_left_out;
wire [0:228] sb_1__1__137_chanx_right_out;
wire [0:228] sb_1__1__137_chany_bottom_out;
wire [0:228] sb_1__1__137_chany_top_out;
wire [0:0] sb_1__1__138_ccff_tail;
wire [0:228] sb_1__1__138_chanx_left_out;
wire [0:228] sb_1__1__138_chanx_right_out;
wire [0:228] sb_1__1__138_chany_bottom_out;
wire [0:228] sb_1__1__138_chany_top_out;
wire [0:0] sb_1__1__139_ccff_tail;
wire [0:228] sb_1__1__139_chanx_left_out;
wire [0:228] sb_1__1__139_chanx_right_out;
wire [0:228] sb_1__1__139_chany_bottom_out;
wire [0:228] sb_1__1__139_chany_top_out;
wire [0:0] sb_1__1__13_ccff_tail;
wire [0:228] sb_1__1__13_chanx_left_out;
wire [0:228] sb_1__1__13_chanx_right_out;
wire [0:228] sb_1__1__13_chany_bottom_out;
wire [0:228] sb_1__1__13_chany_top_out;
wire [0:0] sb_1__1__140_ccff_tail;
wire [0:228] sb_1__1__140_chanx_left_out;
wire [0:228] sb_1__1__140_chanx_right_out;
wire [0:228] sb_1__1__140_chany_bottom_out;
wire [0:228] sb_1__1__140_chany_top_out;
wire [0:0] sb_1__1__141_ccff_tail;
wire [0:228] sb_1__1__141_chanx_left_out;
wire [0:228] sb_1__1__141_chanx_right_out;
wire [0:228] sb_1__1__141_chany_bottom_out;
wire [0:228] sb_1__1__141_chany_top_out;
wire [0:0] sb_1__1__142_ccff_tail;
wire [0:228] sb_1__1__142_chanx_left_out;
wire [0:228] sb_1__1__142_chanx_right_out;
wire [0:228] sb_1__1__142_chany_bottom_out;
wire [0:228] sb_1__1__142_chany_top_out;
wire [0:0] sb_1__1__143_ccff_tail;
wire [0:228] sb_1__1__143_chanx_left_out;
wire [0:228] sb_1__1__143_chanx_right_out;
wire [0:228] sb_1__1__143_chany_bottom_out;
wire [0:228] sb_1__1__143_chany_top_out;
wire [0:0] sb_1__1__144_ccff_tail;
wire [0:228] sb_1__1__144_chanx_left_out;
wire [0:228] sb_1__1__144_chanx_right_out;
wire [0:228] sb_1__1__144_chany_bottom_out;
wire [0:228] sb_1__1__144_chany_top_out;
wire [0:0] sb_1__1__145_ccff_tail;
wire [0:228] sb_1__1__145_chanx_left_out;
wire [0:228] sb_1__1__145_chanx_right_out;
wire [0:228] sb_1__1__145_chany_bottom_out;
wire [0:228] sb_1__1__145_chany_top_out;
wire [0:0] sb_1__1__146_ccff_tail;
wire [0:228] sb_1__1__146_chanx_left_out;
wire [0:228] sb_1__1__146_chanx_right_out;
wire [0:228] sb_1__1__146_chany_bottom_out;
wire [0:228] sb_1__1__146_chany_top_out;
wire [0:0] sb_1__1__147_ccff_tail;
wire [0:228] sb_1__1__147_chanx_left_out;
wire [0:228] sb_1__1__147_chanx_right_out;
wire [0:228] sb_1__1__147_chany_bottom_out;
wire [0:228] sb_1__1__147_chany_top_out;
wire [0:0] sb_1__1__148_ccff_tail;
wire [0:228] sb_1__1__148_chanx_left_out;
wire [0:228] sb_1__1__148_chanx_right_out;
wire [0:228] sb_1__1__148_chany_bottom_out;
wire [0:228] sb_1__1__148_chany_top_out;
wire [0:0] sb_1__1__149_ccff_tail;
wire [0:228] sb_1__1__149_chanx_left_out;
wire [0:228] sb_1__1__149_chanx_right_out;
wire [0:228] sb_1__1__149_chany_bottom_out;
wire [0:228] sb_1__1__149_chany_top_out;
wire [0:0] sb_1__1__14_ccff_tail;
wire [0:228] sb_1__1__14_chanx_left_out;
wire [0:228] sb_1__1__14_chanx_right_out;
wire [0:228] sb_1__1__14_chany_bottom_out;
wire [0:228] sb_1__1__14_chany_top_out;
wire [0:0] sb_1__1__150_ccff_tail;
wire [0:228] sb_1__1__150_chanx_left_out;
wire [0:228] sb_1__1__150_chanx_right_out;
wire [0:228] sb_1__1__150_chany_bottom_out;
wire [0:228] sb_1__1__150_chany_top_out;
wire [0:0] sb_1__1__151_ccff_tail;
wire [0:228] sb_1__1__151_chanx_left_out;
wire [0:228] sb_1__1__151_chanx_right_out;
wire [0:228] sb_1__1__151_chany_bottom_out;
wire [0:228] sb_1__1__151_chany_top_out;
wire [0:0] sb_1__1__152_ccff_tail;
wire [0:228] sb_1__1__152_chanx_left_out;
wire [0:228] sb_1__1__152_chanx_right_out;
wire [0:228] sb_1__1__152_chany_bottom_out;
wire [0:228] sb_1__1__152_chany_top_out;
wire [0:0] sb_1__1__153_ccff_tail;
wire [0:228] sb_1__1__153_chanx_left_out;
wire [0:228] sb_1__1__153_chanx_right_out;
wire [0:228] sb_1__1__153_chany_bottom_out;
wire [0:228] sb_1__1__153_chany_top_out;
wire [0:0] sb_1__1__154_ccff_tail;
wire [0:228] sb_1__1__154_chanx_left_out;
wire [0:228] sb_1__1__154_chanx_right_out;
wire [0:228] sb_1__1__154_chany_bottom_out;
wire [0:228] sb_1__1__154_chany_top_out;
wire [0:0] sb_1__1__155_ccff_tail;
wire [0:228] sb_1__1__155_chanx_left_out;
wire [0:228] sb_1__1__155_chanx_right_out;
wire [0:228] sb_1__1__155_chany_bottom_out;
wire [0:228] sb_1__1__155_chany_top_out;
wire [0:0] sb_1__1__156_ccff_tail;
wire [0:228] sb_1__1__156_chanx_left_out;
wire [0:228] sb_1__1__156_chanx_right_out;
wire [0:228] sb_1__1__156_chany_bottom_out;
wire [0:228] sb_1__1__156_chany_top_out;
wire [0:0] sb_1__1__157_ccff_tail;
wire [0:228] sb_1__1__157_chanx_left_out;
wire [0:228] sb_1__1__157_chanx_right_out;
wire [0:228] sb_1__1__157_chany_bottom_out;
wire [0:228] sb_1__1__157_chany_top_out;
wire [0:0] sb_1__1__158_ccff_tail;
wire [0:228] sb_1__1__158_chanx_left_out;
wire [0:228] sb_1__1__158_chanx_right_out;
wire [0:228] sb_1__1__158_chany_bottom_out;
wire [0:228] sb_1__1__158_chany_top_out;
wire [0:0] sb_1__1__159_ccff_tail;
wire [0:228] sb_1__1__159_chanx_left_out;
wire [0:228] sb_1__1__159_chanx_right_out;
wire [0:228] sb_1__1__159_chany_bottom_out;
wire [0:228] sb_1__1__159_chany_top_out;
wire [0:0] sb_1__1__15_ccff_tail;
wire [0:228] sb_1__1__15_chanx_left_out;
wire [0:228] sb_1__1__15_chanx_right_out;
wire [0:228] sb_1__1__15_chany_bottom_out;
wire [0:228] sb_1__1__15_chany_top_out;
wire [0:0] sb_1__1__160_ccff_tail;
wire [0:228] sb_1__1__160_chanx_left_out;
wire [0:228] sb_1__1__160_chanx_right_out;
wire [0:228] sb_1__1__160_chany_bottom_out;
wire [0:228] sb_1__1__160_chany_top_out;
wire [0:0] sb_1__1__161_ccff_tail;
wire [0:228] sb_1__1__161_chanx_left_out;
wire [0:228] sb_1__1__161_chanx_right_out;
wire [0:228] sb_1__1__161_chany_bottom_out;
wire [0:228] sb_1__1__161_chany_top_out;
wire [0:0] sb_1__1__162_ccff_tail;
wire [0:228] sb_1__1__162_chanx_left_out;
wire [0:228] sb_1__1__162_chanx_right_out;
wire [0:228] sb_1__1__162_chany_bottom_out;
wire [0:228] sb_1__1__162_chany_top_out;
wire [0:0] sb_1__1__163_ccff_tail;
wire [0:228] sb_1__1__163_chanx_left_out;
wire [0:228] sb_1__1__163_chanx_right_out;
wire [0:228] sb_1__1__163_chany_bottom_out;
wire [0:228] sb_1__1__163_chany_top_out;
wire [0:0] sb_1__1__164_ccff_tail;
wire [0:228] sb_1__1__164_chanx_left_out;
wire [0:228] sb_1__1__164_chanx_right_out;
wire [0:228] sb_1__1__164_chany_bottom_out;
wire [0:228] sb_1__1__164_chany_top_out;
wire [0:0] sb_1__1__165_ccff_tail;
wire [0:228] sb_1__1__165_chanx_left_out;
wire [0:228] sb_1__1__165_chanx_right_out;
wire [0:228] sb_1__1__165_chany_bottom_out;
wire [0:228] sb_1__1__165_chany_top_out;
wire [0:0] sb_1__1__166_ccff_tail;
wire [0:228] sb_1__1__166_chanx_left_out;
wire [0:228] sb_1__1__166_chanx_right_out;
wire [0:228] sb_1__1__166_chany_bottom_out;
wire [0:228] sb_1__1__166_chany_top_out;
wire [0:0] sb_1__1__167_ccff_tail;
wire [0:228] sb_1__1__167_chanx_left_out;
wire [0:228] sb_1__1__167_chanx_right_out;
wire [0:228] sb_1__1__167_chany_bottom_out;
wire [0:228] sb_1__1__167_chany_top_out;
wire [0:0] sb_1__1__168_ccff_tail;
wire [0:228] sb_1__1__168_chanx_left_out;
wire [0:228] sb_1__1__168_chanx_right_out;
wire [0:228] sb_1__1__168_chany_bottom_out;
wire [0:228] sb_1__1__168_chany_top_out;
wire [0:0] sb_1__1__169_ccff_tail;
wire [0:228] sb_1__1__169_chanx_left_out;
wire [0:228] sb_1__1__169_chanx_right_out;
wire [0:228] sb_1__1__169_chany_bottom_out;
wire [0:228] sb_1__1__169_chany_top_out;
wire [0:0] sb_1__1__16_ccff_tail;
wire [0:228] sb_1__1__16_chanx_left_out;
wire [0:228] sb_1__1__16_chanx_right_out;
wire [0:228] sb_1__1__16_chany_bottom_out;
wire [0:228] sb_1__1__16_chany_top_out;
wire [0:0] sb_1__1__170_ccff_tail;
wire [0:228] sb_1__1__170_chanx_left_out;
wire [0:228] sb_1__1__170_chanx_right_out;
wire [0:228] sb_1__1__170_chany_bottom_out;
wire [0:228] sb_1__1__170_chany_top_out;
wire [0:0] sb_1__1__171_ccff_tail;
wire [0:228] sb_1__1__171_chanx_left_out;
wire [0:228] sb_1__1__171_chanx_right_out;
wire [0:228] sb_1__1__171_chany_bottom_out;
wire [0:228] sb_1__1__171_chany_top_out;
wire [0:0] sb_1__1__172_ccff_tail;
wire [0:228] sb_1__1__172_chanx_left_out;
wire [0:228] sb_1__1__172_chanx_right_out;
wire [0:228] sb_1__1__172_chany_bottom_out;
wire [0:228] sb_1__1__172_chany_top_out;
wire [0:0] sb_1__1__173_ccff_tail;
wire [0:228] sb_1__1__173_chanx_left_out;
wire [0:228] sb_1__1__173_chanx_right_out;
wire [0:228] sb_1__1__173_chany_bottom_out;
wire [0:228] sb_1__1__173_chany_top_out;
wire [0:0] sb_1__1__174_ccff_tail;
wire [0:228] sb_1__1__174_chanx_left_out;
wire [0:228] sb_1__1__174_chanx_right_out;
wire [0:228] sb_1__1__174_chany_bottom_out;
wire [0:228] sb_1__1__174_chany_top_out;
wire [0:0] sb_1__1__175_ccff_tail;
wire [0:228] sb_1__1__175_chanx_left_out;
wire [0:228] sb_1__1__175_chanx_right_out;
wire [0:228] sb_1__1__175_chany_bottom_out;
wire [0:228] sb_1__1__175_chany_top_out;
wire [0:0] sb_1__1__176_ccff_tail;
wire [0:228] sb_1__1__176_chanx_left_out;
wire [0:228] sb_1__1__176_chanx_right_out;
wire [0:228] sb_1__1__176_chany_bottom_out;
wire [0:228] sb_1__1__176_chany_top_out;
wire [0:0] sb_1__1__177_ccff_tail;
wire [0:228] sb_1__1__177_chanx_left_out;
wire [0:228] sb_1__1__177_chanx_right_out;
wire [0:228] sb_1__1__177_chany_bottom_out;
wire [0:228] sb_1__1__177_chany_top_out;
wire [0:0] sb_1__1__178_ccff_tail;
wire [0:228] sb_1__1__178_chanx_left_out;
wire [0:228] sb_1__1__178_chanx_right_out;
wire [0:228] sb_1__1__178_chany_bottom_out;
wire [0:228] sb_1__1__178_chany_top_out;
wire [0:0] sb_1__1__179_ccff_tail;
wire [0:228] sb_1__1__179_chanx_left_out;
wire [0:228] sb_1__1__179_chanx_right_out;
wire [0:228] sb_1__1__179_chany_bottom_out;
wire [0:228] sb_1__1__179_chany_top_out;
wire [0:0] sb_1__1__17_ccff_tail;
wire [0:228] sb_1__1__17_chanx_left_out;
wire [0:228] sb_1__1__17_chanx_right_out;
wire [0:228] sb_1__1__17_chany_bottom_out;
wire [0:228] sb_1__1__17_chany_top_out;
wire [0:0] sb_1__1__180_ccff_tail;
wire [0:228] sb_1__1__180_chanx_left_out;
wire [0:228] sb_1__1__180_chanx_right_out;
wire [0:228] sb_1__1__180_chany_bottom_out;
wire [0:228] sb_1__1__180_chany_top_out;
wire [0:0] sb_1__1__181_ccff_tail;
wire [0:228] sb_1__1__181_chanx_left_out;
wire [0:228] sb_1__1__181_chanx_right_out;
wire [0:228] sb_1__1__181_chany_bottom_out;
wire [0:228] sb_1__1__181_chany_top_out;
wire [0:0] sb_1__1__182_ccff_tail;
wire [0:228] sb_1__1__182_chanx_left_out;
wire [0:228] sb_1__1__182_chanx_right_out;
wire [0:228] sb_1__1__182_chany_bottom_out;
wire [0:228] sb_1__1__182_chany_top_out;
wire [0:0] sb_1__1__183_ccff_tail;
wire [0:228] sb_1__1__183_chanx_left_out;
wire [0:228] sb_1__1__183_chanx_right_out;
wire [0:228] sb_1__1__183_chany_bottom_out;
wire [0:228] sb_1__1__183_chany_top_out;
wire [0:0] sb_1__1__184_ccff_tail;
wire [0:228] sb_1__1__184_chanx_left_out;
wire [0:228] sb_1__1__184_chanx_right_out;
wire [0:228] sb_1__1__184_chany_bottom_out;
wire [0:228] sb_1__1__184_chany_top_out;
wire [0:0] sb_1__1__185_ccff_tail;
wire [0:228] sb_1__1__185_chanx_left_out;
wire [0:228] sb_1__1__185_chanx_right_out;
wire [0:228] sb_1__1__185_chany_bottom_out;
wire [0:228] sb_1__1__185_chany_top_out;
wire [0:0] sb_1__1__186_ccff_tail;
wire [0:228] sb_1__1__186_chanx_left_out;
wire [0:228] sb_1__1__186_chanx_right_out;
wire [0:228] sb_1__1__186_chany_bottom_out;
wire [0:228] sb_1__1__186_chany_top_out;
wire [0:0] sb_1__1__187_ccff_tail;
wire [0:228] sb_1__1__187_chanx_left_out;
wire [0:228] sb_1__1__187_chanx_right_out;
wire [0:228] sb_1__1__187_chany_bottom_out;
wire [0:228] sb_1__1__187_chany_top_out;
wire [0:0] sb_1__1__188_ccff_tail;
wire [0:228] sb_1__1__188_chanx_left_out;
wire [0:228] sb_1__1__188_chanx_right_out;
wire [0:228] sb_1__1__188_chany_bottom_out;
wire [0:228] sb_1__1__188_chany_top_out;
wire [0:0] sb_1__1__189_ccff_tail;
wire [0:228] sb_1__1__189_chanx_left_out;
wire [0:228] sb_1__1__189_chanx_right_out;
wire [0:228] sb_1__1__189_chany_bottom_out;
wire [0:228] sb_1__1__189_chany_top_out;
wire [0:228] sb_1__1__18_chanx_left_out;
wire [0:228] sb_1__1__18_chanx_right_out;
wire [0:228] sb_1__1__18_chany_bottom_out;
wire [0:228] sb_1__1__18_chany_top_out;
wire [0:0] sb_1__1__190_ccff_tail;
wire [0:228] sb_1__1__190_chanx_left_out;
wire [0:228] sb_1__1__190_chanx_right_out;
wire [0:228] sb_1__1__190_chany_bottom_out;
wire [0:228] sb_1__1__190_chany_top_out;
wire [0:0] sb_1__1__191_ccff_tail;
wire [0:228] sb_1__1__191_chanx_left_out;
wire [0:228] sb_1__1__191_chanx_right_out;
wire [0:228] sb_1__1__191_chany_bottom_out;
wire [0:228] sb_1__1__191_chany_top_out;
wire [0:0] sb_1__1__192_ccff_tail;
wire [0:228] sb_1__1__192_chanx_left_out;
wire [0:228] sb_1__1__192_chanx_right_out;
wire [0:228] sb_1__1__192_chany_bottom_out;
wire [0:228] sb_1__1__192_chany_top_out;
wire [0:0] sb_1__1__193_ccff_tail;
wire [0:228] sb_1__1__193_chanx_left_out;
wire [0:228] sb_1__1__193_chanx_right_out;
wire [0:228] sb_1__1__193_chany_bottom_out;
wire [0:228] sb_1__1__193_chany_top_out;
wire [0:0] sb_1__1__194_ccff_tail;
wire [0:228] sb_1__1__194_chanx_left_out;
wire [0:228] sb_1__1__194_chanx_right_out;
wire [0:228] sb_1__1__194_chany_bottom_out;
wire [0:228] sb_1__1__194_chany_top_out;
wire [0:0] sb_1__1__195_ccff_tail;
wire [0:228] sb_1__1__195_chanx_left_out;
wire [0:228] sb_1__1__195_chanx_right_out;
wire [0:228] sb_1__1__195_chany_bottom_out;
wire [0:228] sb_1__1__195_chany_top_out;
wire [0:0] sb_1__1__196_ccff_tail;
wire [0:228] sb_1__1__196_chanx_left_out;
wire [0:228] sb_1__1__196_chanx_right_out;
wire [0:228] sb_1__1__196_chany_bottom_out;
wire [0:228] sb_1__1__196_chany_top_out;
wire [0:0] sb_1__1__197_ccff_tail;
wire [0:228] sb_1__1__197_chanx_left_out;
wire [0:228] sb_1__1__197_chanx_right_out;
wire [0:228] sb_1__1__197_chany_bottom_out;
wire [0:228] sb_1__1__197_chany_top_out;
wire [0:0] sb_1__1__198_ccff_tail;
wire [0:228] sb_1__1__198_chanx_left_out;
wire [0:228] sb_1__1__198_chanx_right_out;
wire [0:228] sb_1__1__198_chany_bottom_out;
wire [0:228] sb_1__1__198_chany_top_out;
wire [0:0] sb_1__1__199_ccff_tail;
wire [0:228] sb_1__1__199_chanx_left_out;
wire [0:228] sb_1__1__199_chanx_right_out;
wire [0:228] sb_1__1__199_chany_bottom_out;
wire [0:228] sb_1__1__199_chany_top_out;
wire [0:0] sb_1__1__19_ccff_tail;
wire [0:228] sb_1__1__19_chanx_left_out;
wire [0:228] sb_1__1__19_chanx_right_out;
wire [0:228] sb_1__1__19_chany_bottom_out;
wire [0:228] sb_1__1__19_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:228] sb_1__1__1_chanx_left_out;
wire [0:228] sb_1__1__1_chanx_right_out;
wire [0:228] sb_1__1__1_chany_bottom_out;
wire [0:228] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__200_ccff_tail;
wire [0:228] sb_1__1__200_chanx_left_out;
wire [0:228] sb_1__1__200_chanx_right_out;
wire [0:228] sb_1__1__200_chany_bottom_out;
wire [0:228] sb_1__1__200_chany_top_out;
wire [0:0] sb_1__1__201_ccff_tail;
wire [0:228] sb_1__1__201_chanx_left_out;
wire [0:228] sb_1__1__201_chanx_right_out;
wire [0:228] sb_1__1__201_chany_bottom_out;
wire [0:228] sb_1__1__201_chany_top_out;
wire [0:0] sb_1__1__202_ccff_tail;
wire [0:228] sb_1__1__202_chanx_left_out;
wire [0:228] sb_1__1__202_chanx_right_out;
wire [0:228] sb_1__1__202_chany_bottom_out;
wire [0:228] sb_1__1__202_chany_top_out;
wire [0:0] sb_1__1__203_ccff_tail;
wire [0:228] sb_1__1__203_chanx_left_out;
wire [0:228] sb_1__1__203_chanx_right_out;
wire [0:228] sb_1__1__203_chany_bottom_out;
wire [0:228] sb_1__1__203_chany_top_out;
wire [0:0] sb_1__1__204_ccff_tail;
wire [0:228] sb_1__1__204_chanx_left_out;
wire [0:228] sb_1__1__204_chanx_right_out;
wire [0:228] sb_1__1__204_chany_bottom_out;
wire [0:228] sb_1__1__204_chany_top_out;
wire [0:0] sb_1__1__205_ccff_tail;
wire [0:228] sb_1__1__205_chanx_left_out;
wire [0:228] sb_1__1__205_chanx_right_out;
wire [0:228] sb_1__1__205_chany_bottom_out;
wire [0:228] sb_1__1__205_chany_top_out;
wire [0:0] sb_1__1__206_ccff_tail;
wire [0:228] sb_1__1__206_chanx_left_out;
wire [0:228] sb_1__1__206_chanx_right_out;
wire [0:228] sb_1__1__206_chany_bottom_out;
wire [0:228] sb_1__1__206_chany_top_out;
wire [0:0] sb_1__1__207_ccff_tail;
wire [0:228] sb_1__1__207_chanx_left_out;
wire [0:228] sb_1__1__207_chanx_right_out;
wire [0:228] sb_1__1__207_chany_bottom_out;
wire [0:228] sb_1__1__207_chany_top_out;
wire [0:0] sb_1__1__208_ccff_tail;
wire [0:228] sb_1__1__208_chanx_left_out;
wire [0:228] sb_1__1__208_chanx_right_out;
wire [0:228] sb_1__1__208_chany_bottom_out;
wire [0:228] sb_1__1__208_chany_top_out;
wire [0:0] sb_1__1__209_ccff_tail;
wire [0:228] sb_1__1__209_chanx_left_out;
wire [0:228] sb_1__1__209_chanx_right_out;
wire [0:228] sb_1__1__209_chany_bottom_out;
wire [0:228] sb_1__1__209_chany_top_out;
wire [0:0] sb_1__1__20_ccff_tail;
wire [0:228] sb_1__1__20_chanx_left_out;
wire [0:228] sb_1__1__20_chanx_right_out;
wire [0:228] sb_1__1__20_chany_bottom_out;
wire [0:228] sb_1__1__20_chany_top_out;
wire [0:0] sb_1__1__210_ccff_tail;
wire [0:228] sb_1__1__210_chanx_left_out;
wire [0:228] sb_1__1__210_chanx_right_out;
wire [0:228] sb_1__1__210_chany_bottom_out;
wire [0:228] sb_1__1__210_chany_top_out;
wire [0:0] sb_1__1__211_ccff_tail;
wire [0:228] sb_1__1__211_chanx_left_out;
wire [0:228] sb_1__1__211_chanx_right_out;
wire [0:228] sb_1__1__211_chany_bottom_out;
wire [0:228] sb_1__1__211_chany_top_out;
wire [0:0] sb_1__1__212_ccff_tail;
wire [0:228] sb_1__1__212_chanx_left_out;
wire [0:228] sb_1__1__212_chanx_right_out;
wire [0:228] sb_1__1__212_chany_bottom_out;
wire [0:228] sb_1__1__212_chany_top_out;
wire [0:0] sb_1__1__213_ccff_tail;
wire [0:228] sb_1__1__213_chanx_left_out;
wire [0:228] sb_1__1__213_chanx_right_out;
wire [0:228] sb_1__1__213_chany_bottom_out;
wire [0:228] sb_1__1__213_chany_top_out;
wire [0:0] sb_1__1__214_ccff_tail;
wire [0:228] sb_1__1__214_chanx_left_out;
wire [0:228] sb_1__1__214_chanx_right_out;
wire [0:228] sb_1__1__214_chany_bottom_out;
wire [0:228] sb_1__1__214_chany_top_out;
wire [0:0] sb_1__1__215_ccff_tail;
wire [0:228] sb_1__1__215_chanx_left_out;
wire [0:228] sb_1__1__215_chanx_right_out;
wire [0:228] sb_1__1__215_chany_bottom_out;
wire [0:228] sb_1__1__215_chany_top_out;
wire [0:0] sb_1__1__216_ccff_tail;
wire [0:228] sb_1__1__216_chanx_left_out;
wire [0:228] sb_1__1__216_chanx_right_out;
wire [0:228] sb_1__1__216_chany_bottom_out;
wire [0:228] sb_1__1__216_chany_top_out;
wire [0:0] sb_1__1__217_ccff_tail;
wire [0:228] sb_1__1__217_chanx_left_out;
wire [0:228] sb_1__1__217_chanx_right_out;
wire [0:228] sb_1__1__217_chany_bottom_out;
wire [0:228] sb_1__1__217_chany_top_out;
wire [0:0] sb_1__1__218_ccff_tail;
wire [0:228] sb_1__1__218_chanx_left_out;
wire [0:228] sb_1__1__218_chanx_right_out;
wire [0:228] sb_1__1__218_chany_bottom_out;
wire [0:228] sb_1__1__218_chany_top_out;
wire [0:0] sb_1__1__219_ccff_tail;
wire [0:228] sb_1__1__219_chanx_left_out;
wire [0:228] sb_1__1__219_chanx_right_out;
wire [0:228] sb_1__1__219_chany_bottom_out;
wire [0:228] sb_1__1__219_chany_top_out;
wire [0:0] sb_1__1__21_ccff_tail;
wire [0:228] sb_1__1__21_chanx_left_out;
wire [0:228] sb_1__1__21_chanx_right_out;
wire [0:228] sb_1__1__21_chany_bottom_out;
wire [0:228] sb_1__1__21_chany_top_out;
wire [0:0] sb_1__1__220_ccff_tail;
wire [0:228] sb_1__1__220_chanx_left_out;
wire [0:228] sb_1__1__220_chanx_right_out;
wire [0:228] sb_1__1__220_chany_bottom_out;
wire [0:228] sb_1__1__220_chany_top_out;
wire [0:0] sb_1__1__221_ccff_tail;
wire [0:228] sb_1__1__221_chanx_left_out;
wire [0:228] sb_1__1__221_chanx_right_out;
wire [0:228] sb_1__1__221_chany_bottom_out;
wire [0:228] sb_1__1__221_chany_top_out;
wire [0:0] sb_1__1__222_ccff_tail;
wire [0:228] sb_1__1__222_chanx_left_out;
wire [0:228] sb_1__1__222_chanx_right_out;
wire [0:228] sb_1__1__222_chany_bottom_out;
wire [0:228] sb_1__1__222_chany_top_out;
wire [0:0] sb_1__1__223_ccff_tail;
wire [0:228] sb_1__1__223_chanx_left_out;
wire [0:228] sb_1__1__223_chanx_right_out;
wire [0:228] sb_1__1__223_chany_bottom_out;
wire [0:228] sb_1__1__223_chany_top_out;
wire [0:0] sb_1__1__224_ccff_tail;
wire [0:228] sb_1__1__224_chanx_left_out;
wire [0:228] sb_1__1__224_chanx_right_out;
wire [0:228] sb_1__1__224_chany_bottom_out;
wire [0:228] sb_1__1__224_chany_top_out;
wire [0:0] sb_1__1__225_ccff_tail;
wire [0:228] sb_1__1__225_chanx_left_out;
wire [0:228] sb_1__1__225_chanx_right_out;
wire [0:228] sb_1__1__225_chany_bottom_out;
wire [0:228] sb_1__1__225_chany_top_out;
wire [0:0] sb_1__1__226_ccff_tail;
wire [0:228] sb_1__1__226_chanx_left_out;
wire [0:228] sb_1__1__226_chanx_right_out;
wire [0:228] sb_1__1__226_chany_bottom_out;
wire [0:228] sb_1__1__226_chany_top_out;
wire [0:0] sb_1__1__227_ccff_tail;
wire [0:228] sb_1__1__227_chanx_left_out;
wire [0:228] sb_1__1__227_chanx_right_out;
wire [0:228] sb_1__1__227_chany_bottom_out;
wire [0:228] sb_1__1__227_chany_top_out;
wire [0:0] sb_1__1__228_ccff_tail;
wire [0:228] sb_1__1__228_chanx_left_out;
wire [0:228] sb_1__1__228_chanx_right_out;
wire [0:228] sb_1__1__228_chany_bottom_out;
wire [0:228] sb_1__1__228_chany_top_out;
wire [0:0] sb_1__1__229_ccff_tail;
wire [0:228] sb_1__1__229_chanx_left_out;
wire [0:228] sb_1__1__229_chanx_right_out;
wire [0:228] sb_1__1__229_chany_bottom_out;
wire [0:228] sb_1__1__229_chany_top_out;
wire [0:0] sb_1__1__22_ccff_tail;
wire [0:228] sb_1__1__22_chanx_left_out;
wire [0:228] sb_1__1__22_chanx_right_out;
wire [0:228] sb_1__1__22_chany_bottom_out;
wire [0:228] sb_1__1__22_chany_top_out;
wire [0:0] sb_1__1__230_ccff_tail;
wire [0:228] sb_1__1__230_chanx_left_out;
wire [0:228] sb_1__1__230_chanx_right_out;
wire [0:228] sb_1__1__230_chany_bottom_out;
wire [0:228] sb_1__1__230_chany_top_out;
wire [0:0] sb_1__1__231_ccff_tail;
wire [0:228] sb_1__1__231_chanx_left_out;
wire [0:228] sb_1__1__231_chanx_right_out;
wire [0:228] sb_1__1__231_chany_bottom_out;
wire [0:228] sb_1__1__231_chany_top_out;
wire [0:0] sb_1__1__232_ccff_tail;
wire [0:228] sb_1__1__232_chanx_left_out;
wire [0:228] sb_1__1__232_chanx_right_out;
wire [0:228] sb_1__1__232_chany_bottom_out;
wire [0:228] sb_1__1__232_chany_top_out;
wire [0:0] sb_1__1__233_ccff_tail;
wire [0:228] sb_1__1__233_chanx_left_out;
wire [0:228] sb_1__1__233_chanx_right_out;
wire [0:228] sb_1__1__233_chany_bottom_out;
wire [0:228] sb_1__1__233_chany_top_out;
wire [0:0] sb_1__1__234_ccff_tail;
wire [0:228] sb_1__1__234_chanx_left_out;
wire [0:228] sb_1__1__234_chanx_right_out;
wire [0:228] sb_1__1__234_chany_bottom_out;
wire [0:228] sb_1__1__234_chany_top_out;
wire [0:0] sb_1__1__235_ccff_tail;
wire [0:228] sb_1__1__235_chanx_left_out;
wire [0:228] sb_1__1__235_chanx_right_out;
wire [0:228] sb_1__1__235_chany_bottom_out;
wire [0:228] sb_1__1__235_chany_top_out;
wire [0:0] sb_1__1__236_ccff_tail;
wire [0:228] sb_1__1__236_chanx_left_out;
wire [0:228] sb_1__1__236_chanx_right_out;
wire [0:228] sb_1__1__236_chany_bottom_out;
wire [0:228] sb_1__1__236_chany_top_out;
wire [0:0] sb_1__1__237_ccff_tail;
wire [0:228] sb_1__1__237_chanx_left_out;
wire [0:228] sb_1__1__237_chanx_right_out;
wire [0:228] sb_1__1__237_chany_bottom_out;
wire [0:228] sb_1__1__237_chany_top_out;
wire [0:0] sb_1__1__238_ccff_tail;
wire [0:228] sb_1__1__238_chanx_left_out;
wire [0:228] sb_1__1__238_chanx_right_out;
wire [0:228] sb_1__1__238_chany_bottom_out;
wire [0:228] sb_1__1__238_chany_top_out;
wire [0:0] sb_1__1__239_ccff_tail;
wire [0:228] sb_1__1__239_chanx_left_out;
wire [0:228] sb_1__1__239_chanx_right_out;
wire [0:228] sb_1__1__239_chany_bottom_out;
wire [0:228] sb_1__1__239_chany_top_out;
wire [0:0] sb_1__1__23_ccff_tail;
wire [0:228] sb_1__1__23_chanx_left_out;
wire [0:228] sb_1__1__23_chanx_right_out;
wire [0:228] sb_1__1__23_chany_bottom_out;
wire [0:228] sb_1__1__23_chany_top_out;
wire [0:0] sb_1__1__240_ccff_tail;
wire [0:228] sb_1__1__240_chanx_left_out;
wire [0:228] sb_1__1__240_chanx_right_out;
wire [0:228] sb_1__1__240_chany_bottom_out;
wire [0:228] sb_1__1__240_chany_top_out;
wire [0:0] sb_1__1__241_ccff_tail;
wire [0:228] sb_1__1__241_chanx_left_out;
wire [0:228] sb_1__1__241_chanx_right_out;
wire [0:228] sb_1__1__241_chany_bottom_out;
wire [0:228] sb_1__1__241_chany_top_out;
wire [0:0] sb_1__1__242_ccff_tail;
wire [0:228] sb_1__1__242_chanx_left_out;
wire [0:228] sb_1__1__242_chanx_right_out;
wire [0:228] sb_1__1__242_chany_bottom_out;
wire [0:228] sb_1__1__242_chany_top_out;
wire [0:0] sb_1__1__243_ccff_tail;
wire [0:228] sb_1__1__243_chanx_left_out;
wire [0:228] sb_1__1__243_chanx_right_out;
wire [0:228] sb_1__1__243_chany_bottom_out;
wire [0:228] sb_1__1__243_chany_top_out;
wire [0:0] sb_1__1__244_ccff_tail;
wire [0:228] sb_1__1__244_chanx_left_out;
wire [0:228] sb_1__1__244_chanx_right_out;
wire [0:228] sb_1__1__244_chany_bottom_out;
wire [0:228] sb_1__1__244_chany_top_out;
wire [0:0] sb_1__1__245_ccff_tail;
wire [0:228] sb_1__1__245_chanx_left_out;
wire [0:228] sb_1__1__245_chanx_right_out;
wire [0:228] sb_1__1__245_chany_bottom_out;
wire [0:228] sb_1__1__245_chany_top_out;
wire [0:0] sb_1__1__246_ccff_tail;
wire [0:228] sb_1__1__246_chanx_left_out;
wire [0:228] sb_1__1__246_chanx_right_out;
wire [0:228] sb_1__1__246_chany_bottom_out;
wire [0:228] sb_1__1__246_chany_top_out;
wire [0:0] sb_1__1__247_ccff_tail;
wire [0:228] sb_1__1__247_chanx_left_out;
wire [0:228] sb_1__1__247_chanx_right_out;
wire [0:228] sb_1__1__247_chany_bottom_out;
wire [0:228] sb_1__1__247_chany_top_out;
wire [0:0] sb_1__1__248_ccff_tail;
wire [0:228] sb_1__1__248_chanx_left_out;
wire [0:228] sb_1__1__248_chanx_right_out;
wire [0:228] sb_1__1__248_chany_bottom_out;
wire [0:228] sb_1__1__248_chany_top_out;
wire [0:0] sb_1__1__249_ccff_tail;
wire [0:228] sb_1__1__249_chanx_left_out;
wire [0:228] sb_1__1__249_chanx_right_out;
wire [0:228] sb_1__1__249_chany_bottom_out;
wire [0:228] sb_1__1__249_chany_top_out;
wire [0:0] sb_1__1__24_ccff_tail;
wire [0:228] sb_1__1__24_chanx_left_out;
wire [0:228] sb_1__1__24_chanx_right_out;
wire [0:228] sb_1__1__24_chany_bottom_out;
wire [0:228] sb_1__1__24_chany_top_out;
wire [0:0] sb_1__1__250_ccff_tail;
wire [0:228] sb_1__1__250_chanx_left_out;
wire [0:228] sb_1__1__250_chanx_right_out;
wire [0:228] sb_1__1__250_chany_bottom_out;
wire [0:228] sb_1__1__250_chany_top_out;
wire [0:0] sb_1__1__251_ccff_tail;
wire [0:228] sb_1__1__251_chanx_left_out;
wire [0:228] sb_1__1__251_chanx_right_out;
wire [0:228] sb_1__1__251_chany_bottom_out;
wire [0:228] sb_1__1__251_chany_top_out;
wire [0:0] sb_1__1__252_ccff_tail;
wire [0:228] sb_1__1__252_chanx_left_out;
wire [0:228] sb_1__1__252_chanx_right_out;
wire [0:228] sb_1__1__252_chany_bottom_out;
wire [0:228] sb_1__1__252_chany_top_out;
wire [0:0] sb_1__1__253_ccff_tail;
wire [0:228] sb_1__1__253_chanx_left_out;
wire [0:228] sb_1__1__253_chanx_right_out;
wire [0:228] sb_1__1__253_chany_bottom_out;
wire [0:228] sb_1__1__253_chany_top_out;
wire [0:0] sb_1__1__254_ccff_tail;
wire [0:228] sb_1__1__254_chanx_left_out;
wire [0:228] sb_1__1__254_chanx_right_out;
wire [0:228] sb_1__1__254_chany_bottom_out;
wire [0:228] sb_1__1__254_chany_top_out;
wire [0:0] sb_1__1__255_ccff_tail;
wire [0:228] sb_1__1__255_chanx_left_out;
wire [0:228] sb_1__1__255_chanx_right_out;
wire [0:228] sb_1__1__255_chany_bottom_out;
wire [0:228] sb_1__1__255_chany_top_out;
wire [0:0] sb_1__1__256_ccff_tail;
wire [0:228] sb_1__1__256_chanx_left_out;
wire [0:228] sb_1__1__256_chanx_right_out;
wire [0:228] sb_1__1__256_chany_bottom_out;
wire [0:228] sb_1__1__256_chany_top_out;
wire [0:0] sb_1__1__257_ccff_tail;
wire [0:228] sb_1__1__257_chanx_left_out;
wire [0:228] sb_1__1__257_chanx_right_out;
wire [0:228] sb_1__1__257_chany_bottom_out;
wire [0:228] sb_1__1__257_chany_top_out;
wire [0:0] sb_1__1__258_ccff_tail;
wire [0:228] sb_1__1__258_chanx_left_out;
wire [0:228] sb_1__1__258_chanx_right_out;
wire [0:228] sb_1__1__258_chany_bottom_out;
wire [0:228] sb_1__1__258_chany_top_out;
wire [0:0] sb_1__1__259_ccff_tail;
wire [0:228] sb_1__1__259_chanx_left_out;
wire [0:228] sb_1__1__259_chanx_right_out;
wire [0:228] sb_1__1__259_chany_bottom_out;
wire [0:228] sb_1__1__259_chany_top_out;
wire [0:0] sb_1__1__25_ccff_tail;
wire [0:228] sb_1__1__25_chanx_left_out;
wire [0:228] sb_1__1__25_chanx_right_out;
wire [0:228] sb_1__1__25_chany_bottom_out;
wire [0:228] sb_1__1__25_chany_top_out;
wire [0:0] sb_1__1__260_ccff_tail;
wire [0:228] sb_1__1__260_chanx_left_out;
wire [0:228] sb_1__1__260_chanx_right_out;
wire [0:228] sb_1__1__260_chany_bottom_out;
wire [0:228] sb_1__1__260_chany_top_out;
wire [0:0] sb_1__1__261_ccff_tail;
wire [0:228] sb_1__1__261_chanx_left_out;
wire [0:228] sb_1__1__261_chanx_right_out;
wire [0:228] sb_1__1__261_chany_bottom_out;
wire [0:228] sb_1__1__261_chany_top_out;
wire [0:0] sb_1__1__262_ccff_tail;
wire [0:228] sb_1__1__262_chanx_left_out;
wire [0:228] sb_1__1__262_chanx_right_out;
wire [0:228] sb_1__1__262_chany_bottom_out;
wire [0:228] sb_1__1__262_chany_top_out;
wire [0:0] sb_1__1__263_ccff_tail;
wire [0:228] sb_1__1__263_chanx_left_out;
wire [0:228] sb_1__1__263_chanx_right_out;
wire [0:228] sb_1__1__263_chany_bottom_out;
wire [0:228] sb_1__1__263_chany_top_out;
wire [0:0] sb_1__1__264_ccff_tail;
wire [0:228] sb_1__1__264_chanx_left_out;
wire [0:228] sb_1__1__264_chanx_right_out;
wire [0:228] sb_1__1__264_chany_bottom_out;
wire [0:228] sb_1__1__264_chany_top_out;
wire [0:0] sb_1__1__265_ccff_tail;
wire [0:228] sb_1__1__265_chanx_left_out;
wire [0:228] sb_1__1__265_chanx_right_out;
wire [0:228] sb_1__1__265_chany_bottom_out;
wire [0:228] sb_1__1__265_chany_top_out;
wire [0:0] sb_1__1__266_ccff_tail;
wire [0:228] sb_1__1__266_chanx_left_out;
wire [0:228] sb_1__1__266_chanx_right_out;
wire [0:228] sb_1__1__266_chany_bottom_out;
wire [0:228] sb_1__1__266_chany_top_out;
wire [0:0] sb_1__1__267_ccff_tail;
wire [0:228] sb_1__1__267_chanx_left_out;
wire [0:228] sb_1__1__267_chanx_right_out;
wire [0:228] sb_1__1__267_chany_bottom_out;
wire [0:228] sb_1__1__267_chany_top_out;
wire [0:0] sb_1__1__268_ccff_tail;
wire [0:228] sb_1__1__268_chanx_left_out;
wire [0:228] sb_1__1__268_chanx_right_out;
wire [0:228] sb_1__1__268_chany_bottom_out;
wire [0:228] sb_1__1__268_chany_top_out;
wire [0:0] sb_1__1__269_ccff_tail;
wire [0:228] sb_1__1__269_chanx_left_out;
wire [0:228] sb_1__1__269_chanx_right_out;
wire [0:228] sb_1__1__269_chany_bottom_out;
wire [0:228] sb_1__1__269_chany_top_out;
wire [0:0] sb_1__1__26_ccff_tail;
wire [0:228] sb_1__1__26_chanx_left_out;
wire [0:228] sb_1__1__26_chanx_right_out;
wire [0:228] sb_1__1__26_chany_bottom_out;
wire [0:228] sb_1__1__26_chany_top_out;
wire [0:0] sb_1__1__270_ccff_tail;
wire [0:228] sb_1__1__270_chanx_left_out;
wire [0:228] sb_1__1__270_chanx_right_out;
wire [0:228] sb_1__1__270_chany_bottom_out;
wire [0:228] sb_1__1__270_chany_top_out;
wire [0:0] sb_1__1__271_ccff_tail;
wire [0:228] sb_1__1__271_chanx_left_out;
wire [0:228] sb_1__1__271_chanx_right_out;
wire [0:228] sb_1__1__271_chany_bottom_out;
wire [0:228] sb_1__1__271_chany_top_out;
wire [0:0] sb_1__1__272_ccff_tail;
wire [0:228] sb_1__1__272_chanx_left_out;
wire [0:228] sb_1__1__272_chanx_right_out;
wire [0:228] sb_1__1__272_chany_bottom_out;
wire [0:228] sb_1__1__272_chany_top_out;
wire [0:0] sb_1__1__273_ccff_tail;
wire [0:228] sb_1__1__273_chanx_left_out;
wire [0:228] sb_1__1__273_chanx_right_out;
wire [0:228] sb_1__1__273_chany_bottom_out;
wire [0:228] sb_1__1__273_chany_top_out;
wire [0:0] sb_1__1__274_ccff_tail;
wire [0:228] sb_1__1__274_chanx_left_out;
wire [0:228] sb_1__1__274_chanx_right_out;
wire [0:228] sb_1__1__274_chany_bottom_out;
wire [0:228] sb_1__1__274_chany_top_out;
wire [0:0] sb_1__1__275_ccff_tail;
wire [0:228] sb_1__1__275_chanx_left_out;
wire [0:228] sb_1__1__275_chanx_right_out;
wire [0:228] sb_1__1__275_chany_bottom_out;
wire [0:228] sb_1__1__275_chany_top_out;
wire [0:0] sb_1__1__276_ccff_tail;
wire [0:228] sb_1__1__276_chanx_left_out;
wire [0:228] sb_1__1__276_chanx_right_out;
wire [0:228] sb_1__1__276_chany_bottom_out;
wire [0:228] sb_1__1__276_chany_top_out;
wire [0:0] sb_1__1__277_ccff_tail;
wire [0:228] sb_1__1__277_chanx_left_out;
wire [0:228] sb_1__1__277_chanx_right_out;
wire [0:228] sb_1__1__277_chany_bottom_out;
wire [0:228] sb_1__1__277_chany_top_out;
wire [0:0] sb_1__1__278_ccff_tail;
wire [0:228] sb_1__1__278_chanx_left_out;
wire [0:228] sb_1__1__278_chanx_right_out;
wire [0:228] sb_1__1__278_chany_bottom_out;
wire [0:228] sb_1__1__278_chany_top_out;
wire [0:0] sb_1__1__279_ccff_tail;
wire [0:228] sb_1__1__279_chanx_left_out;
wire [0:228] sb_1__1__279_chanx_right_out;
wire [0:228] sb_1__1__279_chany_bottom_out;
wire [0:228] sb_1__1__279_chany_top_out;
wire [0:0] sb_1__1__27_ccff_tail;
wire [0:228] sb_1__1__27_chanx_left_out;
wire [0:228] sb_1__1__27_chanx_right_out;
wire [0:228] sb_1__1__27_chany_bottom_out;
wire [0:228] sb_1__1__27_chany_top_out;
wire [0:0] sb_1__1__280_ccff_tail;
wire [0:228] sb_1__1__280_chanx_left_out;
wire [0:228] sb_1__1__280_chanx_right_out;
wire [0:228] sb_1__1__280_chany_bottom_out;
wire [0:228] sb_1__1__280_chany_top_out;
wire [0:0] sb_1__1__281_ccff_tail;
wire [0:228] sb_1__1__281_chanx_left_out;
wire [0:228] sb_1__1__281_chanx_right_out;
wire [0:228] sb_1__1__281_chany_bottom_out;
wire [0:228] sb_1__1__281_chany_top_out;
wire [0:0] sb_1__1__282_ccff_tail;
wire [0:228] sb_1__1__282_chanx_left_out;
wire [0:228] sb_1__1__282_chanx_right_out;
wire [0:228] sb_1__1__282_chany_bottom_out;
wire [0:228] sb_1__1__282_chany_top_out;
wire [0:0] sb_1__1__283_ccff_tail;
wire [0:228] sb_1__1__283_chanx_left_out;
wire [0:228] sb_1__1__283_chanx_right_out;
wire [0:228] sb_1__1__283_chany_bottom_out;
wire [0:228] sb_1__1__283_chany_top_out;
wire [0:0] sb_1__1__284_ccff_tail;
wire [0:228] sb_1__1__284_chanx_left_out;
wire [0:228] sb_1__1__284_chanx_right_out;
wire [0:228] sb_1__1__284_chany_bottom_out;
wire [0:228] sb_1__1__284_chany_top_out;
wire [0:0] sb_1__1__285_ccff_tail;
wire [0:228] sb_1__1__285_chanx_left_out;
wire [0:228] sb_1__1__285_chanx_right_out;
wire [0:228] sb_1__1__285_chany_bottom_out;
wire [0:228] sb_1__1__285_chany_top_out;
wire [0:0] sb_1__1__286_ccff_tail;
wire [0:228] sb_1__1__286_chanx_left_out;
wire [0:228] sb_1__1__286_chanx_right_out;
wire [0:228] sb_1__1__286_chany_bottom_out;
wire [0:228] sb_1__1__286_chany_top_out;
wire [0:0] sb_1__1__287_ccff_tail;
wire [0:228] sb_1__1__287_chanx_left_out;
wire [0:228] sb_1__1__287_chanx_right_out;
wire [0:228] sb_1__1__287_chany_bottom_out;
wire [0:228] sb_1__1__287_chany_top_out;
wire [0:0] sb_1__1__288_ccff_tail;
wire [0:228] sb_1__1__288_chanx_left_out;
wire [0:228] sb_1__1__288_chanx_right_out;
wire [0:228] sb_1__1__288_chany_bottom_out;
wire [0:228] sb_1__1__288_chany_top_out;
wire [0:0] sb_1__1__289_ccff_tail;
wire [0:228] sb_1__1__289_chanx_left_out;
wire [0:228] sb_1__1__289_chanx_right_out;
wire [0:228] sb_1__1__289_chany_bottom_out;
wire [0:228] sb_1__1__289_chany_top_out;
wire [0:0] sb_1__1__28_ccff_tail;
wire [0:228] sb_1__1__28_chanx_left_out;
wire [0:228] sb_1__1__28_chanx_right_out;
wire [0:228] sb_1__1__28_chany_bottom_out;
wire [0:228] sb_1__1__28_chany_top_out;
wire [0:0] sb_1__1__290_ccff_tail;
wire [0:228] sb_1__1__290_chanx_left_out;
wire [0:228] sb_1__1__290_chanx_right_out;
wire [0:228] sb_1__1__290_chany_bottom_out;
wire [0:228] sb_1__1__290_chany_top_out;
wire [0:0] sb_1__1__291_ccff_tail;
wire [0:228] sb_1__1__291_chanx_left_out;
wire [0:228] sb_1__1__291_chanx_right_out;
wire [0:228] sb_1__1__291_chany_bottom_out;
wire [0:228] sb_1__1__291_chany_top_out;
wire [0:0] sb_1__1__292_ccff_tail;
wire [0:228] sb_1__1__292_chanx_left_out;
wire [0:228] sb_1__1__292_chanx_right_out;
wire [0:228] sb_1__1__292_chany_bottom_out;
wire [0:228] sb_1__1__292_chany_top_out;
wire [0:0] sb_1__1__293_ccff_tail;
wire [0:228] sb_1__1__293_chanx_left_out;
wire [0:228] sb_1__1__293_chanx_right_out;
wire [0:228] sb_1__1__293_chany_bottom_out;
wire [0:228] sb_1__1__293_chany_top_out;
wire [0:0] sb_1__1__294_ccff_tail;
wire [0:228] sb_1__1__294_chanx_left_out;
wire [0:228] sb_1__1__294_chanx_right_out;
wire [0:228] sb_1__1__294_chany_bottom_out;
wire [0:228] sb_1__1__294_chany_top_out;
wire [0:0] sb_1__1__295_ccff_tail;
wire [0:228] sb_1__1__295_chanx_left_out;
wire [0:228] sb_1__1__295_chanx_right_out;
wire [0:228] sb_1__1__295_chany_bottom_out;
wire [0:228] sb_1__1__295_chany_top_out;
wire [0:0] sb_1__1__296_ccff_tail;
wire [0:228] sb_1__1__296_chanx_left_out;
wire [0:228] sb_1__1__296_chanx_right_out;
wire [0:228] sb_1__1__296_chany_bottom_out;
wire [0:228] sb_1__1__296_chany_top_out;
wire [0:0] sb_1__1__297_ccff_tail;
wire [0:228] sb_1__1__297_chanx_left_out;
wire [0:228] sb_1__1__297_chanx_right_out;
wire [0:228] sb_1__1__297_chany_bottom_out;
wire [0:228] sb_1__1__297_chany_top_out;
wire [0:0] sb_1__1__298_ccff_tail;
wire [0:228] sb_1__1__298_chanx_left_out;
wire [0:228] sb_1__1__298_chanx_right_out;
wire [0:228] sb_1__1__298_chany_bottom_out;
wire [0:228] sb_1__1__298_chany_top_out;
wire [0:0] sb_1__1__299_ccff_tail;
wire [0:228] sb_1__1__299_chanx_left_out;
wire [0:228] sb_1__1__299_chanx_right_out;
wire [0:228] sb_1__1__299_chany_bottom_out;
wire [0:228] sb_1__1__299_chany_top_out;
wire [0:0] sb_1__1__29_ccff_tail;
wire [0:228] sb_1__1__29_chanx_left_out;
wire [0:228] sb_1__1__29_chanx_right_out;
wire [0:228] sb_1__1__29_chany_bottom_out;
wire [0:228] sb_1__1__29_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:228] sb_1__1__2_chanx_left_out;
wire [0:228] sb_1__1__2_chanx_right_out;
wire [0:228] sb_1__1__2_chany_bottom_out;
wire [0:228] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__300_ccff_tail;
wire [0:228] sb_1__1__300_chanx_left_out;
wire [0:228] sb_1__1__300_chanx_right_out;
wire [0:228] sb_1__1__300_chany_bottom_out;
wire [0:228] sb_1__1__300_chany_top_out;
wire [0:0] sb_1__1__301_ccff_tail;
wire [0:228] sb_1__1__301_chanx_left_out;
wire [0:228] sb_1__1__301_chanx_right_out;
wire [0:228] sb_1__1__301_chany_bottom_out;
wire [0:228] sb_1__1__301_chany_top_out;
wire [0:0] sb_1__1__302_ccff_tail;
wire [0:228] sb_1__1__302_chanx_left_out;
wire [0:228] sb_1__1__302_chanx_right_out;
wire [0:228] sb_1__1__302_chany_bottom_out;
wire [0:228] sb_1__1__302_chany_top_out;
wire [0:0] sb_1__1__303_ccff_tail;
wire [0:228] sb_1__1__303_chanx_left_out;
wire [0:228] sb_1__1__303_chanx_right_out;
wire [0:228] sb_1__1__303_chany_bottom_out;
wire [0:228] sb_1__1__303_chany_top_out;
wire [0:0] sb_1__1__304_ccff_tail;
wire [0:228] sb_1__1__304_chanx_left_out;
wire [0:228] sb_1__1__304_chanx_right_out;
wire [0:228] sb_1__1__304_chany_bottom_out;
wire [0:228] sb_1__1__304_chany_top_out;
wire [0:0] sb_1__1__305_ccff_tail;
wire [0:228] sb_1__1__305_chanx_left_out;
wire [0:228] sb_1__1__305_chanx_right_out;
wire [0:228] sb_1__1__305_chany_bottom_out;
wire [0:228] sb_1__1__305_chany_top_out;
wire [0:0] sb_1__1__306_ccff_tail;
wire [0:228] sb_1__1__306_chanx_left_out;
wire [0:228] sb_1__1__306_chanx_right_out;
wire [0:228] sb_1__1__306_chany_bottom_out;
wire [0:228] sb_1__1__306_chany_top_out;
wire [0:0] sb_1__1__307_ccff_tail;
wire [0:228] sb_1__1__307_chanx_left_out;
wire [0:228] sb_1__1__307_chanx_right_out;
wire [0:228] sb_1__1__307_chany_bottom_out;
wire [0:228] sb_1__1__307_chany_top_out;
wire [0:0] sb_1__1__308_ccff_tail;
wire [0:228] sb_1__1__308_chanx_left_out;
wire [0:228] sb_1__1__308_chanx_right_out;
wire [0:228] sb_1__1__308_chany_bottom_out;
wire [0:228] sb_1__1__308_chany_top_out;
wire [0:0] sb_1__1__309_ccff_tail;
wire [0:228] sb_1__1__309_chanx_left_out;
wire [0:228] sb_1__1__309_chanx_right_out;
wire [0:228] sb_1__1__309_chany_bottom_out;
wire [0:228] sb_1__1__309_chany_top_out;
wire [0:0] sb_1__1__30_ccff_tail;
wire [0:228] sb_1__1__30_chanx_left_out;
wire [0:228] sb_1__1__30_chanx_right_out;
wire [0:228] sb_1__1__30_chany_bottom_out;
wire [0:228] sb_1__1__30_chany_top_out;
wire [0:0] sb_1__1__310_ccff_tail;
wire [0:228] sb_1__1__310_chanx_left_out;
wire [0:228] sb_1__1__310_chanx_right_out;
wire [0:228] sb_1__1__310_chany_bottom_out;
wire [0:228] sb_1__1__310_chany_top_out;
wire [0:0] sb_1__1__311_ccff_tail;
wire [0:228] sb_1__1__311_chanx_left_out;
wire [0:228] sb_1__1__311_chanx_right_out;
wire [0:228] sb_1__1__311_chany_bottom_out;
wire [0:228] sb_1__1__311_chany_top_out;
wire [0:0] sb_1__1__312_ccff_tail;
wire [0:228] sb_1__1__312_chanx_left_out;
wire [0:228] sb_1__1__312_chanx_right_out;
wire [0:228] sb_1__1__312_chany_bottom_out;
wire [0:228] sb_1__1__312_chany_top_out;
wire [0:0] sb_1__1__313_ccff_tail;
wire [0:228] sb_1__1__313_chanx_left_out;
wire [0:228] sb_1__1__313_chanx_right_out;
wire [0:228] sb_1__1__313_chany_bottom_out;
wire [0:228] sb_1__1__313_chany_top_out;
wire [0:0] sb_1__1__314_ccff_tail;
wire [0:228] sb_1__1__314_chanx_left_out;
wire [0:228] sb_1__1__314_chanx_right_out;
wire [0:228] sb_1__1__314_chany_bottom_out;
wire [0:228] sb_1__1__314_chany_top_out;
wire [0:0] sb_1__1__315_ccff_tail;
wire [0:228] sb_1__1__315_chanx_left_out;
wire [0:228] sb_1__1__315_chanx_right_out;
wire [0:228] sb_1__1__315_chany_bottom_out;
wire [0:228] sb_1__1__315_chany_top_out;
wire [0:0] sb_1__1__316_ccff_tail;
wire [0:228] sb_1__1__316_chanx_left_out;
wire [0:228] sb_1__1__316_chanx_right_out;
wire [0:228] sb_1__1__316_chany_bottom_out;
wire [0:228] sb_1__1__316_chany_top_out;
wire [0:0] sb_1__1__317_ccff_tail;
wire [0:228] sb_1__1__317_chanx_left_out;
wire [0:228] sb_1__1__317_chanx_right_out;
wire [0:228] sb_1__1__317_chany_bottom_out;
wire [0:228] sb_1__1__317_chany_top_out;
wire [0:0] sb_1__1__318_ccff_tail;
wire [0:228] sb_1__1__318_chanx_left_out;
wire [0:228] sb_1__1__318_chanx_right_out;
wire [0:228] sb_1__1__318_chany_bottom_out;
wire [0:228] sb_1__1__318_chany_top_out;
wire [0:0] sb_1__1__319_ccff_tail;
wire [0:228] sb_1__1__319_chanx_left_out;
wire [0:228] sb_1__1__319_chanx_right_out;
wire [0:228] sb_1__1__319_chany_bottom_out;
wire [0:228] sb_1__1__319_chany_top_out;
wire [0:0] sb_1__1__31_ccff_tail;
wire [0:228] sb_1__1__31_chanx_left_out;
wire [0:228] sb_1__1__31_chanx_right_out;
wire [0:228] sb_1__1__31_chany_bottom_out;
wire [0:228] sb_1__1__31_chany_top_out;
wire [0:0] sb_1__1__320_ccff_tail;
wire [0:228] sb_1__1__320_chanx_left_out;
wire [0:228] sb_1__1__320_chanx_right_out;
wire [0:228] sb_1__1__320_chany_bottom_out;
wire [0:228] sb_1__1__320_chany_top_out;
wire [0:0] sb_1__1__321_ccff_tail;
wire [0:228] sb_1__1__321_chanx_left_out;
wire [0:228] sb_1__1__321_chanx_right_out;
wire [0:228] sb_1__1__321_chany_bottom_out;
wire [0:228] sb_1__1__321_chany_top_out;
wire [0:0] sb_1__1__322_ccff_tail;
wire [0:228] sb_1__1__322_chanx_left_out;
wire [0:228] sb_1__1__322_chanx_right_out;
wire [0:228] sb_1__1__322_chany_bottom_out;
wire [0:228] sb_1__1__322_chany_top_out;
wire [0:0] sb_1__1__323_ccff_tail;
wire [0:228] sb_1__1__323_chanx_left_out;
wire [0:228] sb_1__1__323_chanx_right_out;
wire [0:228] sb_1__1__323_chany_bottom_out;
wire [0:228] sb_1__1__323_chany_top_out;
wire [0:0] sb_1__1__324_ccff_tail;
wire [0:228] sb_1__1__324_chanx_left_out;
wire [0:228] sb_1__1__324_chanx_right_out;
wire [0:228] sb_1__1__324_chany_bottom_out;
wire [0:228] sb_1__1__324_chany_top_out;
wire [0:0] sb_1__1__325_ccff_tail;
wire [0:228] sb_1__1__325_chanx_left_out;
wire [0:228] sb_1__1__325_chanx_right_out;
wire [0:228] sb_1__1__325_chany_bottom_out;
wire [0:228] sb_1__1__325_chany_top_out;
wire [0:0] sb_1__1__326_ccff_tail;
wire [0:228] sb_1__1__326_chanx_left_out;
wire [0:228] sb_1__1__326_chanx_right_out;
wire [0:228] sb_1__1__326_chany_bottom_out;
wire [0:228] sb_1__1__326_chany_top_out;
wire [0:0] sb_1__1__327_ccff_tail;
wire [0:228] sb_1__1__327_chanx_left_out;
wire [0:228] sb_1__1__327_chanx_right_out;
wire [0:228] sb_1__1__327_chany_bottom_out;
wire [0:228] sb_1__1__327_chany_top_out;
wire [0:0] sb_1__1__328_ccff_tail;
wire [0:228] sb_1__1__328_chanx_left_out;
wire [0:228] sb_1__1__328_chanx_right_out;
wire [0:228] sb_1__1__328_chany_bottom_out;
wire [0:228] sb_1__1__328_chany_top_out;
wire [0:0] sb_1__1__329_ccff_tail;
wire [0:228] sb_1__1__329_chanx_left_out;
wire [0:228] sb_1__1__329_chanx_right_out;
wire [0:228] sb_1__1__329_chany_bottom_out;
wire [0:228] sb_1__1__329_chany_top_out;
wire [0:0] sb_1__1__32_ccff_tail;
wire [0:228] sb_1__1__32_chanx_left_out;
wire [0:228] sb_1__1__32_chanx_right_out;
wire [0:228] sb_1__1__32_chany_bottom_out;
wire [0:228] sb_1__1__32_chany_top_out;
wire [0:0] sb_1__1__330_ccff_tail;
wire [0:228] sb_1__1__330_chanx_left_out;
wire [0:228] sb_1__1__330_chanx_right_out;
wire [0:228] sb_1__1__330_chany_bottom_out;
wire [0:228] sb_1__1__330_chany_top_out;
wire [0:0] sb_1__1__331_ccff_tail;
wire [0:228] sb_1__1__331_chanx_left_out;
wire [0:228] sb_1__1__331_chanx_right_out;
wire [0:228] sb_1__1__331_chany_bottom_out;
wire [0:228] sb_1__1__331_chany_top_out;
wire [0:0] sb_1__1__332_ccff_tail;
wire [0:228] sb_1__1__332_chanx_left_out;
wire [0:228] sb_1__1__332_chanx_right_out;
wire [0:228] sb_1__1__332_chany_bottom_out;
wire [0:228] sb_1__1__332_chany_top_out;
wire [0:0] sb_1__1__333_ccff_tail;
wire [0:228] sb_1__1__333_chanx_left_out;
wire [0:228] sb_1__1__333_chanx_right_out;
wire [0:228] sb_1__1__333_chany_bottom_out;
wire [0:228] sb_1__1__333_chany_top_out;
wire [0:0] sb_1__1__334_ccff_tail;
wire [0:228] sb_1__1__334_chanx_left_out;
wire [0:228] sb_1__1__334_chanx_right_out;
wire [0:228] sb_1__1__334_chany_bottom_out;
wire [0:228] sb_1__1__334_chany_top_out;
wire [0:0] sb_1__1__335_ccff_tail;
wire [0:228] sb_1__1__335_chanx_left_out;
wire [0:228] sb_1__1__335_chanx_right_out;
wire [0:228] sb_1__1__335_chany_bottom_out;
wire [0:228] sb_1__1__335_chany_top_out;
wire [0:0] sb_1__1__336_ccff_tail;
wire [0:228] sb_1__1__336_chanx_left_out;
wire [0:228] sb_1__1__336_chanx_right_out;
wire [0:228] sb_1__1__336_chany_bottom_out;
wire [0:228] sb_1__1__336_chany_top_out;
wire [0:0] sb_1__1__337_ccff_tail;
wire [0:228] sb_1__1__337_chanx_left_out;
wire [0:228] sb_1__1__337_chanx_right_out;
wire [0:228] sb_1__1__337_chany_bottom_out;
wire [0:228] sb_1__1__337_chany_top_out;
wire [0:0] sb_1__1__338_ccff_tail;
wire [0:228] sb_1__1__338_chanx_left_out;
wire [0:228] sb_1__1__338_chanx_right_out;
wire [0:228] sb_1__1__338_chany_bottom_out;
wire [0:228] sb_1__1__338_chany_top_out;
wire [0:0] sb_1__1__339_ccff_tail;
wire [0:228] sb_1__1__339_chanx_left_out;
wire [0:228] sb_1__1__339_chanx_right_out;
wire [0:228] sb_1__1__339_chany_bottom_out;
wire [0:228] sb_1__1__339_chany_top_out;
wire [0:0] sb_1__1__33_ccff_tail;
wire [0:228] sb_1__1__33_chanx_left_out;
wire [0:228] sb_1__1__33_chanx_right_out;
wire [0:228] sb_1__1__33_chany_bottom_out;
wire [0:228] sb_1__1__33_chany_top_out;
wire [0:0] sb_1__1__340_ccff_tail;
wire [0:228] sb_1__1__340_chanx_left_out;
wire [0:228] sb_1__1__340_chanx_right_out;
wire [0:228] sb_1__1__340_chany_bottom_out;
wire [0:228] sb_1__1__340_chany_top_out;
wire [0:0] sb_1__1__341_ccff_tail;
wire [0:228] sb_1__1__341_chanx_left_out;
wire [0:228] sb_1__1__341_chanx_right_out;
wire [0:228] sb_1__1__341_chany_bottom_out;
wire [0:228] sb_1__1__341_chany_top_out;
wire [0:0] sb_1__1__342_ccff_tail;
wire [0:228] sb_1__1__342_chanx_left_out;
wire [0:228] sb_1__1__342_chanx_right_out;
wire [0:228] sb_1__1__342_chany_bottom_out;
wire [0:228] sb_1__1__342_chany_top_out;
wire [0:0] sb_1__1__343_ccff_tail;
wire [0:228] sb_1__1__343_chanx_left_out;
wire [0:228] sb_1__1__343_chanx_right_out;
wire [0:228] sb_1__1__343_chany_bottom_out;
wire [0:228] sb_1__1__343_chany_top_out;
wire [0:0] sb_1__1__344_ccff_tail;
wire [0:228] sb_1__1__344_chanx_left_out;
wire [0:228] sb_1__1__344_chanx_right_out;
wire [0:228] sb_1__1__344_chany_bottom_out;
wire [0:228] sb_1__1__344_chany_top_out;
wire [0:0] sb_1__1__345_ccff_tail;
wire [0:228] sb_1__1__345_chanx_left_out;
wire [0:228] sb_1__1__345_chanx_right_out;
wire [0:228] sb_1__1__345_chany_bottom_out;
wire [0:228] sb_1__1__345_chany_top_out;
wire [0:0] sb_1__1__346_ccff_tail;
wire [0:228] sb_1__1__346_chanx_left_out;
wire [0:228] sb_1__1__346_chanx_right_out;
wire [0:228] sb_1__1__346_chany_bottom_out;
wire [0:228] sb_1__1__346_chany_top_out;
wire [0:0] sb_1__1__347_ccff_tail;
wire [0:228] sb_1__1__347_chanx_left_out;
wire [0:228] sb_1__1__347_chanx_right_out;
wire [0:228] sb_1__1__347_chany_bottom_out;
wire [0:228] sb_1__1__347_chany_top_out;
wire [0:0] sb_1__1__348_ccff_tail;
wire [0:228] sb_1__1__348_chanx_left_out;
wire [0:228] sb_1__1__348_chanx_right_out;
wire [0:228] sb_1__1__348_chany_bottom_out;
wire [0:228] sb_1__1__348_chany_top_out;
wire [0:0] sb_1__1__349_ccff_tail;
wire [0:228] sb_1__1__349_chanx_left_out;
wire [0:228] sb_1__1__349_chanx_right_out;
wire [0:228] sb_1__1__349_chany_bottom_out;
wire [0:228] sb_1__1__349_chany_top_out;
wire [0:0] sb_1__1__34_ccff_tail;
wire [0:228] sb_1__1__34_chanx_left_out;
wire [0:228] sb_1__1__34_chanx_right_out;
wire [0:228] sb_1__1__34_chany_bottom_out;
wire [0:228] sb_1__1__34_chany_top_out;
wire [0:0] sb_1__1__350_ccff_tail;
wire [0:228] sb_1__1__350_chanx_left_out;
wire [0:228] sb_1__1__350_chanx_right_out;
wire [0:228] sb_1__1__350_chany_bottom_out;
wire [0:228] sb_1__1__350_chany_top_out;
wire [0:0] sb_1__1__351_ccff_tail;
wire [0:228] sb_1__1__351_chanx_left_out;
wire [0:228] sb_1__1__351_chanx_right_out;
wire [0:228] sb_1__1__351_chany_bottom_out;
wire [0:228] sb_1__1__351_chany_top_out;
wire [0:0] sb_1__1__352_ccff_tail;
wire [0:228] sb_1__1__352_chanx_left_out;
wire [0:228] sb_1__1__352_chanx_right_out;
wire [0:228] sb_1__1__352_chany_bottom_out;
wire [0:228] sb_1__1__352_chany_top_out;
wire [0:0] sb_1__1__353_ccff_tail;
wire [0:228] sb_1__1__353_chanx_left_out;
wire [0:228] sb_1__1__353_chanx_right_out;
wire [0:228] sb_1__1__353_chany_bottom_out;
wire [0:228] sb_1__1__353_chany_top_out;
wire [0:0] sb_1__1__354_ccff_tail;
wire [0:228] sb_1__1__354_chanx_left_out;
wire [0:228] sb_1__1__354_chanx_right_out;
wire [0:228] sb_1__1__354_chany_bottom_out;
wire [0:228] sb_1__1__354_chany_top_out;
wire [0:0] sb_1__1__355_ccff_tail;
wire [0:228] sb_1__1__355_chanx_left_out;
wire [0:228] sb_1__1__355_chanx_right_out;
wire [0:228] sb_1__1__355_chany_bottom_out;
wire [0:228] sb_1__1__355_chany_top_out;
wire [0:0] sb_1__1__356_ccff_tail;
wire [0:228] sb_1__1__356_chanx_left_out;
wire [0:228] sb_1__1__356_chanx_right_out;
wire [0:228] sb_1__1__356_chany_bottom_out;
wire [0:228] sb_1__1__356_chany_top_out;
wire [0:0] sb_1__1__357_ccff_tail;
wire [0:228] sb_1__1__357_chanx_left_out;
wire [0:228] sb_1__1__357_chanx_right_out;
wire [0:228] sb_1__1__357_chany_bottom_out;
wire [0:228] sb_1__1__357_chany_top_out;
wire [0:0] sb_1__1__358_ccff_tail;
wire [0:228] sb_1__1__358_chanx_left_out;
wire [0:228] sb_1__1__358_chanx_right_out;
wire [0:228] sb_1__1__358_chany_bottom_out;
wire [0:228] sb_1__1__358_chany_top_out;
wire [0:0] sb_1__1__359_ccff_tail;
wire [0:228] sb_1__1__359_chanx_left_out;
wire [0:228] sb_1__1__359_chanx_right_out;
wire [0:228] sb_1__1__359_chany_bottom_out;
wire [0:228] sb_1__1__359_chany_top_out;
wire [0:0] sb_1__1__35_ccff_tail;
wire [0:228] sb_1__1__35_chanx_left_out;
wire [0:228] sb_1__1__35_chanx_right_out;
wire [0:228] sb_1__1__35_chany_bottom_out;
wire [0:228] sb_1__1__35_chany_top_out;
wire [0:0] sb_1__1__360_ccff_tail;
wire [0:228] sb_1__1__360_chanx_left_out;
wire [0:228] sb_1__1__360_chanx_right_out;
wire [0:228] sb_1__1__360_chany_bottom_out;
wire [0:228] sb_1__1__360_chany_top_out;
wire [0:0] sb_1__1__361_ccff_tail;
wire [0:228] sb_1__1__361_chanx_left_out;
wire [0:228] sb_1__1__361_chanx_right_out;
wire [0:228] sb_1__1__361_chany_bottom_out;
wire [0:228] sb_1__1__361_chany_top_out;
wire [0:0] sb_1__1__362_ccff_tail;
wire [0:228] sb_1__1__362_chanx_left_out;
wire [0:228] sb_1__1__362_chanx_right_out;
wire [0:228] sb_1__1__362_chany_bottom_out;
wire [0:228] sb_1__1__362_chany_top_out;
wire [0:0] sb_1__1__363_ccff_tail;
wire [0:228] sb_1__1__363_chanx_left_out;
wire [0:228] sb_1__1__363_chanx_right_out;
wire [0:228] sb_1__1__363_chany_bottom_out;
wire [0:228] sb_1__1__363_chany_top_out;
wire [0:0] sb_1__1__364_ccff_tail;
wire [0:228] sb_1__1__364_chanx_left_out;
wire [0:228] sb_1__1__364_chanx_right_out;
wire [0:228] sb_1__1__364_chany_bottom_out;
wire [0:228] sb_1__1__364_chany_top_out;
wire [0:0] sb_1__1__365_ccff_tail;
wire [0:228] sb_1__1__365_chanx_left_out;
wire [0:228] sb_1__1__365_chanx_right_out;
wire [0:228] sb_1__1__365_chany_bottom_out;
wire [0:228] sb_1__1__365_chany_top_out;
wire [0:0] sb_1__1__366_ccff_tail;
wire [0:228] sb_1__1__366_chanx_left_out;
wire [0:228] sb_1__1__366_chanx_right_out;
wire [0:228] sb_1__1__366_chany_bottom_out;
wire [0:228] sb_1__1__366_chany_top_out;
wire [0:0] sb_1__1__367_ccff_tail;
wire [0:228] sb_1__1__367_chanx_left_out;
wire [0:228] sb_1__1__367_chanx_right_out;
wire [0:228] sb_1__1__367_chany_bottom_out;
wire [0:228] sb_1__1__367_chany_top_out;
wire [0:0] sb_1__1__368_ccff_tail;
wire [0:228] sb_1__1__368_chanx_left_out;
wire [0:228] sb_1__1__368_chanx_right_out;
wire [0:228] sb_1__1__368_chany_bottom_out;
wire [0:228] sb_1__1__368_chany_top_out;
wire [0:0] sb_1__1__36_ccff_tail;
wire [0:228] sb_1__1__36_chanx_left_out;
wire [0:228] sb_1__1__36_chanx_right_out;
wire [0:228] sb_1__1__36_chany_bottom_out;
wire [0:228] sb_1__1__36_chany_top_out;
wire [0:0] sb_1__1__37_ccff_tail;
wire [0:228] sb_1__1__37_chanx_left_out;
wire [0:228] sb_1__1__37_chanx_right_out;
wire [0:228] sb_1__1__37_chany_bottom_out;
wire [0:228] sb_1__1__37_chany_top_out;
wire [0:0] sb_1__1__38_ccff_tail;
wire [0:228] sb_1__1__38_chanx_left_out;
wire [0:228] sb_1__1__38_chanx_right_out;
wire [0:228] sb_1__1__38_chany_bottom_out;
wire [0:228] sb_1__1__38_chany_top_out;
wire [0:0] sb_1__1__39_ccff_tail;
wire [0:228] sb_1__1__39_chanx_left_out;
wire [0:228] sb_1__1__39_chanx_right_out;
wire [0:228] sb_1__1__39_chany_bottom_out;
wire [0:228] sb_1__1__39_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:228] sb_1__1__3_chanx_left_out;
wire [0:228] sb_1__1__3_chanx_right_out;
wire [0:228] sb_1__1__3_chany_bottom_out;
wire [0:228] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__40_ccff_tail;
wire [0:228] sb_1__1__40_chanx_left_out;
wire [0:228] sb_1__1__40_chanx_right_out;
wire [0:228] sb_1__1__40_chany_bottom_out;
wire [0:228] sb_1__1__40_chany_top_out;
wire [0:0] sb_1__1__41_ccff_tail;
wire [0:228] sb_1__1__41_chanx_left_out;
wire [0:228] sb_1__1__41_chanx_right_out;
wire [0:228] sb_1__1__41_chany_bottom_out;
wire [0:228] sb_1__1__41_chany_top_out;
wire [0:0] sb_1__1__42_ccff_tail;
wire [0:228] sb_1__1__42_chanx_left_out;
wire [0:228] sb_1__1__42_chanx_right_out;
wire [0:228] sb_1__1__42_chany_bottom_out;
wire [0:228] sb_1__1__42_chany_top_out;
wire [0:0] sb_1__1__43_ccff_tail;
wire [0:228] sb_1__1__43_chanx_left_out;
wire [0:228] sb_1__1__43_chanx_right_out;
wire [0:228] sb_1__1__43_chany_bottom_out;
wire [0:228] sb_1__1__43_chany_top_out;
wire [0:0] sb_1__1__44_ccff_tail;
wire [0:228] sb_1__1__44_chanx_left_out;
wire [0:228] sb_1__1__44_chanx_right_out;
wire [0:228] sb_1__1__44_chany_bottom_out;
wire [0:228] sb_1__1__44_chany_top_out;
wire [0:0] sb_1__1__45_ccff_tail;
wire [0:228] sb_1__1__45_chanx_left_out;
wire [0:228] sb_1__1__45_chanx_right_out;
wire [0:228] sb_1__1__45_chany_bottom_out;
wire [0:228] sb_1__1__45_chany_top_out;
wire [0:0] sb_1__1__46_ccff_tail;
wire [0:228] sb_1__1__46_chanx_left_out;
wire [0:228] sb_1__1__46_chanx_right_out;
wire [0:228] sb_1__1__46_chany_bottom_out;
wire [0:228] sb_1__1__46_chany_top_out;
wire [0:0] sb_1__1__47_ccff_tail;
wire [0:228] sb_1__1__47_chanx_left_out;
wire [0:228] sb_1__1__47_chanx_right_out;
wire [0:228] sb_1__1__47_chany_bottom_out;
wire [0:228] sb_1__1__47_chany_top_out;
wire [0:0] sb_1__1__48_ccff_tail;
wire [0:228] sb_1__1__48_chanx_left_out;
wire [0:228] sb_1__1__48_chanx_right_out;
wire [0:228] sb_1__1__48_chany_bottom_out;
wire [0:228] sb_1__1__48_chany_top_out;
wire [0:0] sb_1__1__49_ccff_tail;
wire [0:228] sb_1__1__49_chanx_left_out;
wire [0:228] sb_1__1__49_chanx_right_out;
wire [0:228] sb_1__1__49_chany_bottom_out;
wire [0:228] sb_1__1__49_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:228] sb_1__1__4_chanx_left_out;
wire [0:228] sb_1__1__4_chanx_right_out;
wire [0:228] sb_1__1__4_chany_bottom_out;
wire [0:228] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__50_ccff_tail;
wire [0:228] sb_1__1__50_chanx_left_out;
wire [0:228] sb_1__1__50_chanx_right_out;
wire [0:228] sb_1__1__50_chany_bottom_out;
wire [0:228] sb_1__1__50_chany_top_out;
wire [0:0] sb_1__1__51_ccff_tail;
wire [0:228] sb_1__1__51_chanx_left_out;
wire [0:228] sb_1__1__51_chanx_right_out;
wire [0:228] sb_1__1__51_chany_bottom_out;
wire [0:228] sb_1__1__51_chany_top_out;
wire [0:0] sb_1__1__52_ccff_tail;
wire [0:228] sb_1__1__52_chanx_left_out;
wire [0:228] sb_1__1__52_chanx_right_out;
wire [0:228] sb_1__1__52_chany_bottom_out;
wire [0:228] sb_1__1__52_chany_top_out;
wire [0:0] sb_1__1__53_ccff_tail;
wire [0:228] sb_1__1__53_chanx_left_out;
wire [0:228] sb_1__1__53_chanx_right_out;
wire [0:228] sb_1__1__53_chany_bottom_out;
wire [0:228] sb_1__1__53_chany_top_out;
wire [0:0] sb_1__1__54_ccff_tail;
wire [0:228] sb_1__1__54_chanx_left_out;
wire [0:228] sb_1__1__54_chanx_right_out;
wire [0:228] sb_1__1__54_chany_bottom_out;
wire [0:228] sb_1__1__54_chany_top_out;
wire [0:0] sb_1__1__55_ccff_tail;
wire [0:228] sb_1__1__55_chanx_left_out;
wire [0:228] sb_1__1__55_chanx_right_out;
wire [0:228] sb_1__1__55_chany_bottom_out;
wire [0:228] sb_1__1__55_chany_top_out;
wire [0:0] sb_1__1__56_ccff_tail;
wire [0:228] sb_1__1__56_chanx_left_out;
wire [0:228] sb_1__1__56_chanx_right_out;
wire [0:228] sb_1__1__56_chany_bottom_out;
wire [0:228] sb_1__1__56_chany_top_out;
wire [0:0] sb_1__1__57_ccff_tail;
wire [0:228] sb_1__1__57_chanx_left_out;
wire [0:228] sb_1__1__57_chanx_right_out;
wire [0:228] sb_1__1__57_chany_bottom_out;
wire [0:228] sb_1__1__57_chany_top_out;
wire [0:0] sb_1__1__58_ccff_tail;
wire [0:228] sb_1__1__58_chanx_left_out;
wire [0:228] sb_1__1__58_chanx_right_out;
wire [0:228] sb_1__1__58_chany_bottom_out;
wire [0:228] sb_1__1__58_chany_top_out;
wire [0:0] sb_1__1__59_ccff_tail;
wire [0:228] sb_1__1__59_chanx_left_out;
wire [0:228] sb_1__1__59_chanx_right_out;
wire [0:228] sb_1__1__59_chany_bottom_out;
wire [0:228] sb_1__1__59_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:228] sb_1__1__5_chanx_left_out;
wire [0:228] sb_1__1__5_chanx_right_out;
wire [0:228] sb_1__1__5_chany_bottom_out;
wire [0:228] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__60_ccff_tail;
wire [0:228] sb_1__1__60_chanx_left_out;
wire [0:228] sb_1__1__60_chanx_right_out;
wire [0:228] sb_1__1__60_chany_bottom_out;
wire [0:228] sb_1__1__60_chany_top_out;
wire [0:0] sb_1__1__61_ccff_tail;
wire [0:228] sb_1__1__61_chanx_left_out;
wire [0:228] sb_1__1__61_chanx_right_out;
wire [0:228] sb_1__1__61_chany_bottom_out;
wire [0:228] sb_1__1__61_chany_top_out;
wire [0:0] sb_1__1__62_ccff_tail;
wire [0:228] sb_1__1__62_chanx_left_out;
wire [0:228] sb_1__1__62_chanx_right_out;
wire [0:228] sb_1__1__62_chany_bottom_out;
wire [0:228] sb_1__1__62_chany_top_out;
wire [0:0] sb_1__1__63_ccff_tail;
wire [0:228] sb_1__1__63_chanx_left_out;
wire [0:228] sb_1__1__63_chanx_right_out;
wire [0:228] sb_1__1__63_chany_bottom_out;
wire [0:228] sb_1__1__63_chany_top_out;
wire [0:0] sb_1__1__64_ccff_tail;
wire [0:228] sb_1__1__64_chanx_left_out;
wire [0:228] sb_1__1__64_chanx_right_out;
wire [0:228] sb_1__1__64_chany_bottom_out;
wire [0:228] sb_1__1__64_chany_top_out;
wire [0:0] sb_1__1__65_ccff_tail;
wire [0:228] sb_1__1__65_chanx_left_out;
wire [0:228] sb_1__1__65_chanx_right_out;
wire [0:228] sb_1__1__65_chany_bottom_out;
wire [0:228] sb_1__1__65_chany_top_out;
wire [0:0] sb_1__1__66_ccff_tail;
wire [0:228] sb_1__1__66_chanx_left_out;
wire [0:228] sb_1__1__66_chanx_right_out;
wire [0:228] sb_1__1__66_chany_bottom_out;
wire [0:228] sb_1__1__66_chany_top_out;
wire [0:0] sb_1__1__67_ccff_tail;
wire [0:228] sb_1__1__67_chanx_left_out;
wire [0:228] sb_1__1__67_chanx_right_out;
wire [0:228] sb_1__1__67_chany_bottom_out;
wire [0:228] sb_1__1__67_chany_top_out;
wire [0:0] sb_1__1__68_ccff_tail;
wire [0:228] sb_1__1__68_chanx_left_out;
wire [0:228] sb_1__1__68_chanx_right_out;
wire [0:228] sb_1__1__68_chany_bottom_out;
wire [0:228] sb_1__1__68_chany_top_out;
wire [0:0] sb_1__1__69_ccff_tail;
wire [0:228] sb_1__1__69_chanx_left_out;
wire [0:228] sb_1__1__69_chanx_right_out;
wire [0:228] sb_1__1__69_chany_bottom_out;
wire [0:228] sb_1__1__69_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:228] sb_1__1__6_chanx_left_out;
wire [0:228] sb_1__1__6_chanx_right_out;
wire [0:228] sb_1__1__6_chany_bottom_out;
wire [0:228] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__70_ccff_tail;
wire [0:228] sb_1__1__70_chanx_left_out;
wire [0:228] sb_1__1__70_chanx_right_out;
wire [0:228] sb_1__1__70_chany_bottom_out;
wire [0:228] sb_1__1__70_chany_top_out;
wire [0:0] sb_1__1__71_ccff_tail;
wire [0:228] sb_1__1__71_chanx_left_out;
wire [0:228] sb_1__1__71_chanx_right_out;
wire [0:228] sb_1__1__71_chany_bottom_out;
wire [0:228] sb_1__1__71_chany_top_out;
wire [0:0] sb_1__1__72_ccff_tail;
wire [0:228] sb_1__1__72_chanx_left_out;
wire [0:228] sb_1__1__72_chanx_right_out;
wire [0:228] sb_1__1__72_chany_bottom_out;
wire [0:228] sb_1__1__72_chany_top_out;
wire [0:0] sb_1__1__73_ccff_tail;
wire [0:228] sb_1__1__73_chanx_left_out;
wire [0:228] sb_1__1__73_chanx_right_out;
wire [0:228] sb_1__1__73_chany_bottom_out;
wire [0:228] sb_1__1__73_chany_top_out;
wire [0:0] sb_1__1__74_ccff_tail;
wire [0:228] sb_1__1__74_chanx_left_out;
wire [0:228] sb_1__1__74_chanx_right_out;
wire [0:228] sb_1__1__74_chany_bottom_out;
wire [0:228] sb_1__1__74_chany_top_out;
wire [0:0] sb_1__1__75_ccff_tail;
wire [0:228] sb_1__1__75_chanx_left_out;
wire [0:228] sb_1__1__75_chanx_right_out;
wire [0:228] sb_1__1__75_chany_bottom_out;
wire [0:228] sb_1__1__75_chany_top_out;
wire [0:0] sb_1__1__76_ccff_tail;
wire [0:228] sb_1__1__76_chanx_left_out;
wire [0:228] sb_1__1__76_chanx_right_out;
wire [0:228] sb_1__1__76_chany_bottom_out;
wire [0:228] sb_1__1__76_chany_top_out;
wire [0:0] sb_1__1__77_ccff_tail;
wire [0:228] sb_1__1__77_chanx_left_out;
wire [0:228] sb_1__1__77_chanx_right_out;
wire [0:228] sb_1__1__77_chany_bottom_out;
wire [0:228] sb_1__1__77_chany_top_out;
wire [0:0] sb_1__1__78_ccff_tail;
wire [0:228] sb_1__1__78_chanx_left_out;
wire [0:228] sb_1__1__78_chanx_right_out;
wire [0:228] sb_1__1__78_chany_bottom_out;
wire [0:228] sb_1__1__78_chany_top_out;
wire [0:0] sb_1__1__79_ccff_tail;
wire [0:228] sb_1__1__79_chanx_left_out;
wire [0:228] sb_1__1__79_chanx_right_out;
wire [0:228] sb_1__1__79_chany_bottom_out;
wire [0:228] sb_1__1__79_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:228] sb_1__1__7_chanx_left_out;
wire [0:228] sb_1__1__7_chanx_right_out;
wire [0:228] sb_1__1__7_chany_bottom_out;
wire [0:228] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__80_ccff_tail;
wire [0:228] sb_1__1__80_chanx_left_out;
wire [0:228] sb_1__1__80_chanx_right_out;
wire [0:228] sb_1__1__80_chany_bottom_out;
wire [0:228] sb_1__1__80_chany_top_out;
wire [0:0] sb_1__1__81_ccff_tail;
wire [0:228] sb_1__1__81_chanx_left_out;
wire [0:228] sb_1__1__81_chanx_right_out;
wire [0:228] sb_1__1__81_chany_bottom_out;
wire [0:228] sb_1__1__81_chany_top_out;
wire [0:0] sb_1__1__82_ccff_tail;
wire [0:228] sb_1__1__82_chanx_left_out;
wire [0:228] sb_1__1__82_chanx_right_out;
wire [0:228] sb_1__1__82_chany_bottom_out;
wire [0:228] sb_1__1__82_chany_top_out;
wire [0:0] sb_1__1__83_ccff_tail;
wire [0:228] sb_1__1__83_chanx_left_out;
wire [0:228] sb_1__1__83_chanx_right_out;
wire [0:228] sb_1__1__83_chany_bottom_out;
wire [0:228] sb_1__1__83_chany_top_out;
wire [0:0] sb_1__1__84_ccff_tail;
wire [0:228] sb_1__1__84_chanx_left_out;
wire [0:228] sb_1__1__84_chanx_right_out;
wire [0:228] sb_1__1__84_chany_bottom_out;
wire [0:228] sb_1__1__84_chany_top_out;
wire [0:0] sb_1__1__85_ccff_tail;
wire [0:228] sb_1__1__85_chanx_left_out;
wire [0:228] sb_1__1__85_chanx_right_out;
wire [0:228] sb_1__1__85_chany_bottom_out;
wire [0:228] sb_1__1__85_chany_top_out;
wire [0:0] sb_1__1__86_ccff_tail;
wire [0:228] sb_1__1__86_chanx_left_out;
wire [0:228] sb_1__1__86_chanx_right_out;
wire [0:228] sb_1__1__86_chany_bottom_out;
wire [0:228] sb_1__1__86_chany_top_out;
wire [0:0] sb_1__1__87_ccff_tail;
wire [0:228] sb_1__1__87_chanx_left_out;
wire [0:228] sb_1__1__87_chanx_right_out;
wire [0:228] sb_1__1__87_chany_bottom_out;
wire [0:228] sb_1__1__87_chany_top_out;
wire [0:0] sb_1__1__88_ccff_tail;
wire [0:228] sb_1__1__88_chanx_left_out;
wire [0:228] sb_1__1__88_chanx_right_out;
wire [0:228] sb_1__1__88_chany_bottom_out;
wire [0:228] sb_1__1__88_chany_top_out;
wire [0:0] sb_1__1__89_ccff_tail;
wire [0:228] sb_1__1__89_chanx_left_out;
wire [0:228] sb_1__1__89_chanx_right_out;
wire [0:228] sb_1__1__89_chany_bottom_out;
wire [0:228] sb_1__1__89_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:228] sb_1__1__8_chanx_left_out;
wire [0:228] sb_1__1__8_chanx_right_out;
wire [0:228] sb_1__1__8_chany_bottom_out;
wire [0:228] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__1__90_ccff_tail;
wire [0:228] sb_1__1__90_chanx_left_out;
wire [0:228] sb_1__1__90_chanx_right_out;
wire [0:228] sb_1__1__90_chany_bottom_out;
wire [0:228] sb_1__1__90_chany_top_out;
wire [0:0] sb_1__1__91_ccff_tail;
wire [0:228] sb_1__1__91_chanx_left_out;
wire [0:228] sb_1__1__91_chanx_right_out;
wire [0:228] sb_1__1__91_chany_bottom_out;
wire [0:228] sb_1__1__91_chany_top_out;
wire [0:0] sb_1__1__92_ccff_tail;
wire [0:228] sb_1__1__92_chanx_left_out;
wire [0:228] sb_1__1__92_chanx_right_out;
wire [0:228] sb_1__1__92_chany_bottom_out;
wire [0:228] sb_1__1__92_chany_top_out;
wire [0:0] sb_1__1__93_ccff_tail;
wire [0:228] sb_1__1__93_chanx_left_out;
wire [0:228] sb_1__1__93_chanx_right_out;
wire [0:228] sb_1__1__93_chany_bottom_out;
wire [0:228] sb_1__1__93_chany_top_out;
wire [0:0] sb_1__1__94_ccff_tail;
wire [0:228] sb_1__1__94_chanx_left_out;
wire [0:228] sb_1__1__94_chanx_right_out;
wire [0:228] sb_1__1__94_chany_bottom_out;
wire [0:228] sb_1__1__94_chany_top_out;
wire [0:0] sb_1__1__95_ccff_tail;
wire [0:228] sb_1__1__95_chanx_left_out;
wire [0:228] sb_1__1__95_chanx_right_out;
wire [0:228] sb_1__1__95_chany_bottom_out;
wire [0:228] sb_1__1__95_chany_top_out;
wire [0:0] sb_1__1__96_ccff_tail;
wire [0:228] sb_1__1__96_chanx_left_out;
wire [0:228] sb_1__1__96_chanx_right_out;
wire [0:228] sb_1__1__96_chany_bottom_out;
wire [0:228] sb_1__1__96_chany_top_out;
wire [0:0] sb_1__1__97_ccff_tail;
wire [0:228] sb_1__1__97_chanx_left_out;
wire [0:228] sb_1__1__97_chanx_right_out;
wire [0:228] sb_1__1__97_chany_bottom_out;
wire [0:228] sb_1__1__97_chany_top_out;
wire [0:0] sb_1__1__98_ccff_tail;
wire [0:228] sb_1__1__98_chanx_left_out;
wire [0:228] sb_1__1__98_chanx_right_out;
wire [0:228] sb_1__1__98_chany_bottom_out;
wire [0:228] sb_1__1__98_chany_top_out;
wire [0:0] sb_1__1__99_ccff_tail;
wire [0:228] sb_1__1__99_chanx_left_out;
wire [0:228] sb_1__1__99_chanx_right_out;
wire [0:228] sb_1__1__99_chany_bottom_out;
wire [0:228] sb_1__1__99_chany_top_out;
wire [0:0] sb_1__1__9_ccff_tail;
wire [0:228] sb_1__1__9_chanx_left_out;
wire [0:228] sb_1__1__9_chanx_right_out;
wire [0:228] sb_1__1__9_chany_bottom_out;
wire [0:228] sb_1__1__9_chany_top_out;
wire [0:0] sb_1__22__0_ccff_tail;
wire [0:228] sb_1__22__0_chanx_left_out;
wire [0:228] sb_1__22__0_chanx_right_out;
wire [0:228] sb_1__22__0_chany_bottom_out;
wire [0:0] sb_1__22__10_ccff_tail;
wire [0:228] sb_1__22__10_chanx_left_out;
wire [0:228] sb_1__22__10_chanx_right_out;
wire [0:228] sb_1__22__10_chany_bottom_out;
wire [0:0] sb_1__22__11_ccff_tail;
wire [0:228] sb_1__22__11_chanx_left_out;
wire [0:228] sb_1__22__11_chanx_right_out;
wire [0:228] sb_1__22__11_chany_bottom_out;
wire [0:0] sb_1__22__12_ccff_tail;
wire [0:228] sb_1__22__12_chanx_left_out;
wire [0:228] sb_1__22__12_chanx_right_out;
wire [0:228] sb_1__22__12_chany_bottom_out;
wire [0:0] sb_1__22__13_ccff_tail;
wire [0:228] sb_1__22__13_chanx_left_out;
wire [0:228] sb_1__22__13_chanx_right_out;
wire [0:228] sb_1__22__13_chany_bottom_out;
wire [0:0] sb_1__22__14_ccff_tail;
wire [0:228] sb_1__22__14_chanx_left_out;
wire [0:228] sb_1__22__14_chanx_right_out;
wire [0:228] sb_1__22__14_chany_bottom_out;
wire [0:0] sb_1__22__15_ccff_tail;
wire [0:228] sb_1__22__15_chanx_left_out;
wire [0:228] sb_1__22__15_chanx_right_out;
wire [0:228] sb_1__22__15_chany_bottom_out;
wire [0:0] sb_1__22__16_ccff_tail;
wire [0:228] sb_1__22__16_chanx_left_out;
wire [0:228] sb_1__22__16_chanx_right_out;
wire [0:228] sb_1__22__16_chany_bottom_out;
wire [0:0] sb_1__22__17_ccff_tail;
wire [0:228] sb_1__22__17_chanx_left_out;
wire [0:228] sb_1__22__17_chanx_right_out;
wire [0:228] sb_1__22__17_chany_bottom_out;
wire [0:0] sb_1__22__18_ccff_tail;
wire [0:228] sb_1__22__18_chanx_left_out;
wire [0:228] sb_1__22__18_chanx_right_out;
wire [0:228] sb_1__22__18_chany_bottom_out;
wire [0:0] sb_1__22__19_ccff_tail;
wire [0:228] sb_1__22__19_chanx_left_out;
wire [0:228] sb_1__22__19_chanx_right_out;
wire [0:228] sb_1__22__19_chany_bottom_out;
wire [0:0] sb_1__22__1_ccff_tail;
wire [0:228] sb_1__22__1_chanx_left_out;
wire [0:228] sb_1__22__1_chanx_right_out;
wire [0:228] sb_1__22__1_chany_bottom_out;
wire [0:0] sb_1__22__20_ccff_tail;
wire [0:228] sb_1__22__20_chanx_left_out;
wire [0:228] sb_1__22__20_chanx_right_out;
wire [0:228] sb_1__22__20_chany_bottom_out;
wire [0:0] sb_1__22__2_ccff_tail;
wire [0:228] sb_1__22__2_chanx_left_out;
wire [0:228] sb_1__22__2_chanx_right_out;
wire [0:228] sb_1__22__2_chany_bottom_out;
wire [0:0] sb_1__22__3_ccff_tail;
wire [0:228] sb_1__22__3_chanx_left_out;
wire [0:228] sb_1__22__3_chanx_right_out;
wire [0:228] sb_1__22__3_chany_bottom_out;
wire [0:0] sb_1__22__4_ccff_tail;
wire [0:228] sb_1__22__4_chanx_left_out;
wire [0:228] sb_1__22__4_chanx_right_out;
wire [0:228] sb_1__22__4_chany_bottom_out;
wire [0:0] sb_1__22__5_ccff_tail;
wire [0:228] sb_1__22__5_chanx_left_out;
wire [0:228] sb_1__22__5_chanx_right_out;
wire [0:228] sb_1__22__5_chany_bottom_out;
wire [0:0] sb_1__22__6_ccff_tail;
wire [0:228] sb_1__22__6_chanx_left_out;
wire [0:228] sb_1__22__6_chanx_right_out;
wire [0:228] sb_1__22__6_chany_bottom_out;
wire [0:0] sb_1__22__7_ccff_tail;
wire [0:228] sb_1__22__7_chanx_left_out;
wire [0:228] sb_1__22__7_chanx_right_out;
wire [0:228] sb_1__22__7_chany_bottom_out;
wire [0:0] sb_1__22__8_ccff_tail;
wire [0:228] sb_1__22__8_chanx_left_out;
wire [0:228] sb_1__22__8_chanx_right_out;
wire [0:228] sb_1__22__8_chany_bottom_out;
wire [0:0] sb_1__22__9_ccff_tail;
wire [0:228] sb_1__22__9_chanx_left_out;
wire [0:228] sb_1__22__9_chanx_right_out;
wire [0:228] sb_1__22__9_chany_bottom_out;
wire [0:0] sb_1__4__0_ccff_tail;
wire [0:228] sb_1__4__0_chanx_left_out;
wire [0:228] sb_1__4__0_chanx_right_out;
wire [0:228] sb_1__4__0_chany_bottom_out;
wire [0:228] sb_1__4__0_chany_top_out;
wire [0:0] sb_1__4__10_ccff_tail;
wire [0:228] sb_1__4__10_chanx_left_out;
wire [0:228] sb_1__4__10_chanx_right_out;
wire [0:228] sb_1__4__10_chany_bottom_out;
wire [0:228] sb_1__4__10_chany_top_out;
wire [0:0] sb_1__4__11_ccff_tail;
wire [0:228] sb_1__4__11_chanx_left_out;
wire [0:228] sb_1__4__11_chanx_right_out;
wire [0:228] sb_1__4__11_chany_bottom_out;
wire [0:228] sb_1__4__11_chany_top_out;
wire [0:0] sb_1__4__12_ccff_tail;
wire [0:228] sb_1__4__12_chanx_left_out;
wire [0:228] sb_1__4__12_chanx_right_out;
wire [0:228] sb_1__4__12_chany_bottom_out;
wire [0:228] sb_1__4__12_chany_top_out;
wire [0:0] sb_1__4__13_ccff_tail;
wire [0:228] sb_1__4__13_chanx_left_out;
wire [0:228] sb_1__4__13_chanx_right_out;
wire [0:228] sb_1__4__13_chany_bottom_out;
wire [0:228] sb_1__4__13_chany_top_out;
wire [0:0] sb_1__4__14_ccff_tail;
wire [0:228] sb_1__4__14_chanx_left_out;
wire [0:228] sb_1__4__14_chanx_right_out;
wire [0:228] sb_1__4__14_chany_bottom_out;
wire [0:228] sb_1__4__14_chany_top_out;
wire [0:0] sb_1__4__15_ccff_tail;
wire [0:228] sb_1__4__15_chanx_left_out;
wire [0:228] sb_1__4__15_chanx_right_out;
wire [0:228] sb_1__4__15_chany_bottom_out;
wire [0:228] sb_1__4__15_chany_top_out;
wire [0:0] sb_1__4__16_ccff_tail;
wire [0:228] sb_1__4__16_chanx_left_out;
wire [0:228] sb_1__4__16_chanx_right_out;
wire [0:228] sb_1__4__16_chany_bottom_out;
wire [0:228] sb_1__4__16_chany_top_out;
wire [0:0] sb_1__4__17_ccff_tail;
wire [0:228] sb_1__4__17_chanx_left_out;
wire [0:228] sb_1__4__17_chanx_right_out;
wire [0:228] sb_1__4__17_chany_bottom_out;
wire [0:228] sb_1__4__17_chany_top_out;
wire [0:0] sb_1__4__18_ccff_tail;
wire [0:228] sb_1__4__18_chanx_left_out;
wire [0:228] sb_1__4__18_chanx_right_out;
wire [0:228] sb_1__4__18_chany_bottom_out;
wire [0:228] sb_1__4__18_chany_top_out;
wire [0:0] sb_1__4__19_ccff_tail;
wire [0:228] sb_1__4__19_chanx_left_out;
wire [0:228] sb_1__4__19_chanx_right_out;
wire [0:228] sb_1__4__19_chany_bottom_out;
wire [0:228] sb_1__4__19_chany_top_out;
wire [0:0] sb_1__4__1_ccff_tail;
wire [0:228] sb_1__4__1_chanx_left_out;
wire [0:228] sb_1__4__1_chanx_right_out;
wire [0:228] sb_1__4__1_chany_bottom_out;
wire [0:228] sb_1__4__1_chany_top_out;
wire [0:0] sb_1__4__20_ccff_tail;
wire [0:228] sb_1__4__20_chanx_left_out;
wire [0:228] sb_1__4__20_chanx_right_out;
wire [0:228] sb_1__4__20_chany_bottom_out;
wire [0:228] sb_1__4__20_chany_top_out;
wire [0:0] sb_1__4__2_ccff_tail;
wire [0:228] sb_1__4__2_chanx_left_out;
wire [0:228] sb_1__4__2_chanx_right_out;
wire [0:228] sb_1__4__2_chany_bottom_out;
wire [0:228] sb_1__4__2_chany_top_out;
wire [0:0] sb_1__4__3_ccff_tail;
wire [0:228] sb_1__4__3_chanx_left_out;
wire [0:228] sb_1__4__3_chanx_right_out;
wire [0:228] sb_1__4__3_chany_bottom_out;
wire [0:228] sb_1__4__3_chany_top_out;
wire [0:0] sb_1__4__4_ccff_tail;
wire [0:228] sb_1__4__4_chanx_left_out;
wire [0:228] sb_1__4__4_chanx_right_out;
wire [0:228] sb_1__4__4_chany_bottom_out;
wire [0:228] sb_1__4__4_chany_top_out;
wire [0:0] sb_1__4__5_ccff_tail;
wire [0:228] sb_1__4__5_chanx_left_out;
wire [0:228] sb_1__4__5_chanx_right_out;
wire [0:228] sb_1__4__5_chany_bottom_out;
wire [0:228] sb_1__4__5_chany_top_out;
wire [0:0] sb_1__4__6_ccff_tail;
wire [0:228] sb_1__4__6_chanx_left_out;
wire [0:228] sb_1__4__6_chanx_right_out;
wire [0:228] sb_1__4__6_chany_bottom_out;
wire [0:228] sb_1__4__6_chany_top_out;
wire [0:0] sb_1__4__7_ccff_tail;
wire [0:228] sb_1__4__7_chanx_left_out;
wire [0:228] sb_1__4__7_chanx_right_out;
wire [0:228] sb_1__4__7_chany_bottom_out;
wire [0:228] sb_1__4__7_chany_top_out;
wire [0:0] sb_1__4__8_ccff_tail;
wire [0:228] sb_1__4__8_chanx_left_out;
wire [0:228] sb_1__4__8_chanx_right_out;
wire [0:228] sb_1__4__8_chany_bottom_out;
wire [0:228] sb_1__4__8_chany_top_out;
wire [0:0] sb_1__4__9_ccff_tail;
wire [0:228] sb_1__4__9_chanx_left_out;
wire [0:228] sb_1__4__9_chanx_right_out;
wire [0:228] sb_1__4__9_chany_bottom_out;
wire [0:228] sb_1__4__9_chany_top_out;
wire [0:0] sb_1__5__0_ccff_tail;
wire [0:228] sb_1__5__0_chanx_left_out;
wire [0:228] sb_1__5__0_chanx_right_out;
wire [0:228] sb_1__5__0_chany_bottom_out;
wire [0:228] sb_1__5__0_chany_top_out;
wire [0:0] sb_1__5__10_ccff_tail;
wire [0:228] sb_1__5__10_chanx_left_out;
wire [0:228] sb_1__5__10_chanx_right_out;
wire [0:228] sb_1__5__10_chany_bottom_out;
wire [0:228] sb_1__5__10_chany_top_out;
wire [0:0] sb_1__5__11_ccff_tail;
wire [0:228] sb_1__5__11_chanx_left_out;
wire [0:228] sb_1__5__11_chanx_right_out;
wire [0:228] sb_1__5__11_chany_bottom_out;
wire [0:228] sb_1__5__11_chany_top_out;
wire [0:0] sb_1__5__12_ccff_tail;
wire [0:228] sb_1__5__12_chanx_left_out;
wire [0:228] sb_1__5__12_chanx_right_out;
wire [0:228] sb_1__5__12_chany_bottom_out;
wire [0:228] sb_1__5__12_chany_top_out;
wire [0:0] sb_1__5__13_ccff_tail;
wire [0:228] sb_1__5__13_chanx_left_out;
wire [0:228] sb_1__5__13_chanx_right_out;
wire [0:228] sb_1__5__13_chany_bottom_out;
wire [0:228] sb_1__5__13_chany_top_out;
wire [0:0] sb_1__5__14_ccff_tail;
wire [0:228] sb_1__5__14_chanx_left_out;
wire [0:228] sb_1__5__14_chanx_right_out;
wire [0:228] sb_1__5__14_chany_bottom_out;
wire [0:228] sb_1__5__14_chany_top_out;
wire [0:0] sb_1__5__1_ccff_tail;
wire [0:228] sb_1__5__1_chanx_left_out;
wire [0:228] sb_1__5__1_chanx_right_out;
wire [0:228] sb_1__5__1_chany_bottom_out;
wire [0:228] sb_1__5__1_chany_top_out;
wire [0:0] sb_1__5__2_ccff_tail;
wire [0:228] sb_1__5__2_chanx_left_out;
wire [0:228] sb_1__5__2_chanx_right_out;
wire [0:228] sb_1__5__2_chany_bottom_out;
wire [0:228] sb_1__5__2_chany_top_out;
wire [0:0] sb_1__5__3_ccff_tail;
wire [0:228] sb_1__5__3_chanx_left_out;
wire [0:228] sb_1__5__3_chanx_right_out;
wire [0:228] sb_1__5__3_chany_bottom_out;
wire [0:228] sb_1__5__3_chany_top_out;
wire [0:0] sb_1__5__4_ccff_tail;
wire [0:228] sb_1__5__4_chanx_left_out;
wire [0:228] sb_1__5__4_chanx_right_out;
wire [0:228] sb_1__5__4_chany_bottom_out;
wire [0:228] sb_1__5__4_chany_top_out;
wire [0:0] sb_1__5__5_ccff_tail;
wire [0:228] sb_1__5__5_chanx_left_out;
wire [0:228] sb_1__5__5_chanx_right_out;
wire [0:228] sb_1__5__5_chany_bottom_out;
wire [0:228] sb_1__5__5_chany_top_out;
wire [0:0] sb_1__5__6_ccff_tail;
wire [0:228] sb_1__5__6_chanx_left_out;
wire [0:228] sb_1__5__6_chanx_right_out;
wire [0:228] sb_1__5__6_chany_bottom_out;
wire [0:228] sb_1__5__6_chany_top_out;
wire [0:0] sb_1__5__7_ccff_tail;
wire [0:228] sb_1__5__7_chanx_left_out;
wire [0:228] sb_1__5__7_chanx_right_out;
wire [0:228] sb_1__5__7_chany_bottom_out;
wire [0:228] sb_1__5__7_chany_top_out;
wire [0:0] sb_1__5__8_ccff_tail;
wire [0:228] sb_1__5__8_chanx_left_out;
wire [0:228] sb_1__5__8_chanx_right_out;
wire [0:228] sb_1__5__8_chany_bottom_out;
wire [0:228] sb_1__5__8_chany_top_out;
wire [0:0] sb_1__5__9_ccff_tail;
wire [0:228] sb_1__5__9_chanx_left_out;
wire [0:228] sb_1__5__9_chanx_right_out;
wire [0:228] sb_1__5__9_chany_bottom_out;
wire [0:228] sb_1__5__9_chany_top_out;
wire [0:0] sb_22__0__0_ccff_tail;
wire [0:228] sb_22__0__0_chanx_left_out;
wire [0:228] sb_22__0__0_chany_top_out;
wire [0:0] sb_22__1__0_ccff_tail;
wire [0:228] sb_22__1__0_chanx_left_out;
wire [0:228] sb_22__1__0_chany_bottom_out;
wire [0:228] sb_22__1__0_chany_top_out;
wire [0:0] sb_22__1__10_ccff_tail;
wire [0:228] sb_22__1__10_chanx_left_out;
wire [0:228] sb_22__1__10_chany_bottom_out;
wire [0:228] sb_22__1__10_chany_top_out;
wire [0:0] sb_22__1__11_ccff_tail;
wire [0:228] sb_22__1__11_chanx_left_out;
wire [0:228] sb_22__1__11_chany_bottom_out;
wire [0:228] sb_22__1__11_chany_top_out;
wire [0:0] sb_22__1__12_ccff_tail;
wire [0:228] sb_22__1__12_chanx_left_out;
wire [0:228] sb_22__1__12_chany_bottom_out;
wire [0:228] sb_22__1__12_chany_top_out;
wire [0:0] sb_22__1__13_ccff_tail;
wire [0:228] sb_22__1__13_chanx_left_out;
wire [0:228] sb_22__1__13_chany_bottom_out;
wire [0:228] sb_22__1__13_chany_top_out;
wire [0:0] sb_22__1__14_ccff_tail;
wire [0:228] sb_22__1__14_chanx_left_out;
wire [0:228] sb_22__1__14_chany_bottom_out;
wire [0:228] sb_22__1__14_chany_top_out;
wire [0:0] sb_22__1__15_ccff_tail;
wire [0:228] sb_22__1__15_chanx_left_out;
wire [0:228] sb_22__1__15_chany_bottom_out;
wire [0:228] sb_22__1__15_chany_top_out;
wire [0:0] sb_22__1__16_ccff_tail;
wire [0:228] sb_22__1__16_chanx_left_out;
wire [0:228] sb_22__1__16_chany_bottom_out;
wire [0:228] sb_22__1__16_chany_top_out;
wire [0:0] sb_22__1__17_ccff_tail;
wire [0:228] sb_22__1__17_chanx_left_out;
wire [0:228] sb_22__1__17_chany_bottom_out;
wire [0:228] sb_22__1__17_chany_top_out;
wire [0:0] sb_22__1__18_ccff_tail;
wire [0:228] sb_22__1__18_chanx_left_out;
wire [0:228] sb_22__1__18_chany_bottom_out;
wire [0:228] sb_22__1__18_chany_top_out;
wire [0:0] sb_22__1__1_ccff_tail;
wire [0:228] sb_22__1__1_chanx_left_out;
wire [0:228] sb_22__1__1_chany_bottom_out;
wire [0:228] sb_22__1__1_chany_top_out;
wire [0:0] sb_22__1__2_ccff_tail;
wire [0:228] sb_22__1__2_chanx_left_out;
wire [0:228] sb_22__1__2_chany_bottom_out;
wire [0:228] sb_22__1__2_chany_top_out;
wire [0:0] sb_22__1__3_ccff_tail;
wire [0:228] sb_22__1__3_chanx_left_out;
wire [0:228] sb_22__1__3_chany_bottom_out;
wire [0:228] sb_22__1__3_chany_top_out;
wire [0:0] sb_22__1__4_ccff_tail;
wire [0:228] sb_22__1__4_chanx_left_out;
wire [0:228] sb_22__1__4_chany_bottom_out;
wire [0:228] sb_22__1__4_chany_top_out;
wire [0:0] sb_22__1__5_ccff_tail;
wire [0:228] sb_22__1__5_chanx_left_out;
wire [0:228] sb_22__1__5_chany_bottom_out;
wire [0:228] sb_22__1__5_chany_top_out;
wire [0:0] sb_22__1__6_ccff_tail;
wire [0:228] sb_22__1__6_chanx_left_out;
wire [0:228] sb_22__1__6_chany_bottom_out;
wire [0:228] sb_22__1__6_chany_top_out;
wire [0:0] sb_22__1__7_ccff_tail;
wire [0:228] sb_22__1__7_chanx_left_out;
wire [0:228] sb_22__1__7_chany_bottom_out;
wire [0:228] sb_22__1__7_chany_top_out;
wire [0:0] sb_22__1__8_ccff_tail;
wire [0:228] sb_22__1__8_chanx_left_out;
wire [0:228] sb_22__1__8_chany_bottom_out;
wire [0:228] sb_22__1__8_chany_top_out;
wire [0:0] sb_22__1__9_ccff_tail;
wire [0:228] sb_22__1__9_chanx_left_out;
wire [0:228] sb_22__1__9_chany_bottom_out;
wire [0:228] sb_22__1__9_chany_top_out;
wire [0:0] sb_22__22__0_ccff_tail;
wire [0:228] sb_22__22__0_chanx_left_out;
wire [0:228] sb_22__22__0_chany_bottom_out;
wire [0:0] sb_22__4__0_ccff_tail;
wire [0:228] sb_22__4__0_chanx_left_out;
wire [0:228] sb_22__4__0_chany_bottom_out;
wire [0:228] sb_22__4__0_chany_top_out;
wire [0:0] sb_22__5__0_ccff_tail;
wire [0:228] sb_22__5__0_chanx_left_out;
wire [0:228] sb_22__5__0_chany_bottom_out;
wire [0:228] sb_22__5__0_chany_top_out;
wire [0:0] sb_2__2__0_ccff_tail;
wire [0:228] sb_2__2__0_chanx_left_out;
wire [0:228] sb_2__2__0_chanx_right_out;
wire [0:228] sb_2__2__0_chany_bottom_out;
wire [0:228] sb_2__2__0_chany_top_out;
wire [0:0] sb_2__2__1_ccff_tail;
wire [0:228] sb_2__2__1_chanx_left_out;
wire [0:228] sb_2__2__1_chanx_right_out;
wire [0:228] sb_2__2__1_chany_bottom_out;
wire [0:228] sb_2__2__1_chany_top_out;
wire [0:0] sb_2__2__2_ccff_tail;
wire [0:228] sb_2__2__2_chanx_left_out;
wire [0:228] sb_2__2__2_chanx_right_out;
wire [0:228] sb_2__2__2_chany_bottom_out;
wire [0:228] sb_2__2__2_chany_top_out;
wire [0:0] sb_2__2__3_ccff_tail;
wire [0:228] sb_2__2__3_chanx_left_out;
wire [0:228] sb_2__2__3_chanx_right_out;
wire [0:228] sb_2__2__3_chany_bottom_out;
wire [0:228] sb_2__2__3_chany_top_out;
wire [0:0] sb_2__2__4_ccff_tail;
wire [0:228] sb_2__2__4_chanx_left_out;
wire [0:228] sb_2__2__4_chanx_right_out;
wire [0:228] sb_2__2__4_chany_bottom_out;
wire [0:228] sb_2__2__4_chany_top_out;
wire [0:0] sb_2__2__5_ccff_tail;
wire [0:228] sb_2__2__5_chanx_left_out;
wire [0:228] sb_2__2__5_chanx_right_out;
wire [0:228] sb_2__2__5_chany_bottom_out;
wire [0:228] sb_2__2__5_chany_top_out;
wire [0:0] sb_2__3__0_ccff_tail;
wire [0:228] sb_2__3__0_chanx_left_out;
wire [0:228] sb_2__3__0_chanx_right_out;
wire [0:228] sb_2__3__0_chany_bottom_out;
wire [0:228] sb_2__3__0_chany_top_out;
wire [0:0] sb_2__3__1_ccff_tail;
wire [0:228] sb_2__3__1_chanx_left_out;
wire [0:228] sb_2__3__1_chanx_right_out;
wire [0:228] sb_2__3__1_chany_bottom_out;
wire [0:228] sb_2__3__1_chany_top_out;
wire [0:0] sb_2__3__2_ccff_tail;
wire [0:228] sb_2__3__2_chanx_left_out;
wire [0:228] sb_2__3__2_chanx_right_out;
wire [0:228] sb_2__3__2_chany_bottom_out;
wire [0:228] sb_2__3__2_chany_top_out;
wire [0:0] sb_2__3__3_ccff_tail;
wire [0:228] sb_2__3__3_chanx_left_out;
wire [0:228] sb_2__3__3_chanx_right_out;
wire [0:228] sb_2__3__3_chany_bottom_out;
wire [0:228] sb_2__3__3_chany_top_out;
wire [0:0] sb_2__3__4_ccff_tail;
wire [0:228] sb_2__3__4_chanx_left_out;
wire [0:228] sb_2__3__4_chanx_right_out;
wire [0:228] sb_2__3__4_chany_bottom_out;
wire [0:228] sb_2__3__4_chany_top_out;
wire [0:0] sb_2__3__5_ccff_tail;
wire [0:228] sb_2__3__5_chanx_left_out;
wire [0:228] sb_2__3__5_chanx_right_out;
wire [0:228] sb_2__3__5_chany_bottom_out;
wire [0:228] sb_2__3__5_chany_top_out;
wire [0:0] sb_2__3__6_ccff_tail;
wire [0:228] sb_2__3__6_chanx_left_out;
wire [0:228] sb_2__3__6_chanx_right_out;
wire [0:228] sb_2__3__6_chany_bottom_out;
wire [0:228] sb_2__3__6_chany_top_out;
wire [0:0] sb_2__3__7_ccff_tail;
wire [0:228] sb_2__3__7_chanx_left_out;
wire [0:228] sb_2__3__7_chanx_right_out;
wire [0:228] sb_2__3__7_chany_bottom_out;
wire [0:228] sb_2__3__7_chany_top_out;
wire [0:0] sb_2__3__8_ccff_tail;
wire [0:228] sb_2__3__8_chanx_left_out;
wire [0:228] sb_2__3__8_chanx_right_out;
wire [0:228] sb_2__3__8_chany_bottom_out;
wire [0:228] sb_2__3__8_chany_top_out;
wire [0:0] sb_2__5__0_ccff_tail;
wire [0:228] sb_2__5__0_chanx_left_out;
wire [0:228] sb_2__5__0_chanx_right_out;
wire [0:228] sb_2__5__0_chany_bottom_out;
wire [0:228] sb_2__5__0_chany_top_out;
wire [0:0] sb_2__5__1_ccff_tail;
wire [0:228] sb_2__5__1_chanx_left_out;
wire [0:228] sb_2__5__1_chanx_right_out;
wire [0:228] sb_2__5__1_chany_bottom_out;
wire [0:228] sb_2__5__1_chany_top_out;
wire [0:0] sb_2__5__2_ccff_tail;
wire [0:228] sb_2__5__2_chanx_left_out;
wire [0:228] sb_2__5__2_chanx_right_out;
wire [0:228] sb_2__5__2_chany_bottom_out;
wire [0:228] sb_2__5__2_chany_top_out;
wire [0:0] sb_3__2__0_ccff_tail;
wire [0:228] sb_3__2__0_chanx_left_out;
wire [0:228] sb_3__2__0_chanx_right_out;
wire [0:228] sb_3__2__0_chany_bottom_out;
wire [0:228] sb_3__2__0_chany_top_out;
wire [0:0] sb_3__2__1_ccff_tail;
wire [0:228] sb_3__2__1_chanx_left_out;
wire [0:228] sb_3__2__1_chanx_right_out;
wire [0:228] sb_3__2__1_chany_bottom_out;
wire [0:228] sb_3__2__1_chany_top_out;
wire [0:0] sb_3__2__2_ccff_tail;
wire [0:228] sb_3__2__2_chanx_left_out;
wire [0:228] sb_3__2__2_chanx_right_out;
wire [0:228] sb_3__2__2_chany_bottom_out;
wire [0:228] sb_3__2__2_chany_top_out;
wire [0:0] sb_3__2__3_ccff_tail;
wire [0:228] sb_3__2__3_chanx_left_out;
wire [0:228] sb_3__2__3_chanx_right_out;
wire [0:228] sb_3__2__3_chany_bottom_out;
wire [0:228] sb_3__2__3_chany_top_out;
wire [0:0] sb_3__2__4_ccff_tail;
wire [0:228] sb_3__2__4_chanx_left_out;
wire [0:228] sb_3__2__4_chanx_right_out;
wire [0:228] sb_3__2__4_chany_bottom_out;
wire [0:228] sb_3__2__4_chany_top_out;
wire [0:0] sb_3__2__5_ccff_tail;
wire [0:228] sb_3__2__5_chanx_left_out;
wire [0:228] sb_3__2__5_chanx_right_out;
wire [0:228] sb_3__2__5_chany_bottom_out;
wire [0:228] sb_3__2__5_chany_top_out;
wire [0:0] sb_3__3__0_ccff_tail;
wire [0:228] sb_3__3__0_chanx_left_out;
wire [0:228] sb_3__3__0_chanx_right_out;
wire [0:228] sb_3__3__0_chany_bottom_out;
wire [0:228] sb_3__3__0_chany_top_out;
wire [0:0] sb_3__3__1_ccff_tail;
wire [0:228] sb_3__3__1_chanx_left_out;
wire [0:228] sb_3__3__1_chanx_right_out;
wire [0:228] sb_3__3__1_chany_bottom_out;
wire [0:228] sb_3__3__1_chany_top_out;
wire [0:0] sb_3__3__2_ccff_tail;
wire [0:228] sb_3__3__2_chanx_left_out;
wire [0:228] sb_3__3__2_chanx_right_out;
wire [0:228] sb_3__3__2_chany_bottom_out;
wire [0:228] sb_3__3__2_chany_top_out;
wire [0:0] sb_3__3__3_ccff_tail;
wire [0:228] sb_3__3__3_chanx_left_out;
wire [0:228] sb_3__3__3_chanx_right_out;
wire [0:228] sb_3__3__3_chany_bottom_out;
wire [0:228] sb_3__3__3_chany_top_out;
wire [0:0] sb_3__3__4_ccff_tail;
wire [0:228] sb_3__3__4_chanx_left_out;
wire [0:228] sb_3__3__4_chanx_right_out;
wire [0:228] sb_3__3__4_chany_bottom_out;
wire [0:228] sb_3__3__4_chany_top_out;
wire [0:0] sb_3__3__5_ccff_tail;
wire [0:228] sb_3__3__5_chanx_left_out;
wire [0:228] sb_3__3__5_chanx_right_out;
wire [0:228] sb_3__3__5_chany_bottom_out;
wire [0:228] sb_3__3__5_chany_top_out;
wire [0:0] sb_3__3__6_ccff_tail;
wire [0:228] sb_3__3__6_chanx_left_out;
wire [0:228] sb_3__3__6_chanx_right_out;
wire [0:228] sb_3__3__6_chany_bottom_out;
wire [0:228] sb_3__3__6_chany_top_out;
wire [0:0] sb_3__3__7_ccff_tail;
wire [0:228] sb_3__3__7_chanx_left_out;
wire [0:228] sb_3__3__7_chanx_right_out;
wire [0:228] sb_3__3__7_chany_bottom_out;
wire [0:228] sb_3__3__7_chany_top_out;
wire [0:0] sb_3__3__8_ccff_tail;
wire [0:228] sb_3__3__8_chanx_left_out;
wire [0:228] sb_3__3__8_chanx_right_out;
wire [0:228] sb_3__3__8_chany_bottom_out;
wire [0:228] sb_3__3__8_chany_top_out;
wire [0:0] sb_3__5__0_ccff_tail;
wire [0:228] sb_3__5__0_chanx_left_out;
wire [0:228] sb_3__5__0_chanx_right_out;
wire [0:228] sb_3__5__0_chany_bottom_out;
wire [0:228] sb_3__5__0_chany_top_out;
wire [0:0] sb_3__5__1_ccff_tail;
wire [0:228] sb_3__5__1_chanx_left_out;
wire [0:228] sb_3__5__1_chanx_right_out;
wire [0:228] sb_3__5__1_chany_bottom_out;
wire [0:228] sb_3__5__1_chany_top_out;
wire [0:0] sb_3__5__2_ccff_tail;
wire [0:228] sb_3__5__2_chanx_left_out;
wire [0:228] sb_3__5__2_chanx_right_out;
wire [0:228] sb_3__5__2_chany_bottom_out;
wire [0:228] sb_3__5__2_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_4__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_top grid_io_top_5__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_4_ccff_tail));

	grid_io_top grid_io_top_6__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_5_ccff_tail));

	grid_io_top grid_io_top_7__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__6_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_6_ccff_tail));

	grid_io_top grid_io_top_8__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__7_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_7_ccff_tail));

	grid_io_top grid_io_top_9__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__8_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_8_ccff_tail));

	grid_io_top grid_io_top_10__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__9_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_9_ccff_tail));

	grid_io_top grid_io_top_11__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__10_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_10_ccff_tail));

	grid_io_top grid_io_top_12__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__11_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_11_ccff_tail));

	grid_io_top grid_io_top_13__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__12_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_12_ccff_tail));

	grid_io_top grid_io_top_14__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__13_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_13_ccff_tail));

	grid_io_top grid_io_top_15__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__14_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_14_ccff_tail));

	grid_io_top grid_io_top_16__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__15_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_15_ccff_tail));

	grid_io_top grid_io_top_17__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[128:135]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__16_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_16_ccff_tail));

	grid_io_top grid_io_top_18__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[136:143]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__17_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_17_ccff_tail));

	grid_io_top grid_io_top_19__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[144:151]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__18_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_18_ccff_tail));

	grid_io_top grid_io_top_20__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[152:159]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__19_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_19_ccff_tail));

	grid_io_top grid_io_top_21__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[160:167]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__20_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_20_ccff_tail));

	grid_io_top grid_io_top_22__23_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[168:175]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__22__21_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_21_ccff_tail));

	grid_io_right grid_io_right_23__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[176:183]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_23__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[184:191]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_23__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[192:199]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_23__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[200:207]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right grid_io_right_23__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[208:215]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right grid_io_right_23__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[216:223]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_right grid_io_right_23__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[224:231]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_6_ccff_tail));

	grid_io_right grid_io_right_23__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[232:239]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_7_ccff_tail));

	grid_io_right grid_io_right_23__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[240:247]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_9_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8_ccff_tail));

	grid_io_right grid_io_right_23__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[248:255]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_10_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_9_ccff_tail));

	grid_io_right grid_io_right_23__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[256:263]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_11_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_10_ccff_tail));

	grid_io_right grid_io_right_23__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[264:271]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_12_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_11_ccff_tail));

	grid_io_right grid_io_right_23__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[272:279]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_13_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_12_ccff_tail));

	grid_io_right grid_io_right_23__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[280:287]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_14_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_13_ccff_tail));

	grid_io_right grid_io_right_23__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[288:295]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_15_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_14_ccff_tail));

	grid_io_right grid_io_right_23__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[296:303]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_16_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_15_ccff_tail));

	grid_io_right grid_io_right_23__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[304:311]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_17_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_16_ccff_tail));

	grid_io_right grid_io_right_23__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[312:319]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_18_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_17_ccff_tail));

	grid_io_right grid_io_right_23__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[320:327]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_19_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_18_ccff_tail));

	grid_io_right grid_io_right_23__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[328:335]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_20_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_19_ccff_tail));

	grid_io_right grid_io_right_23__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[336:343]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_21_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_20_ccff_tail));

	grid_io_right grid_io_right_23__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[344:351]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_21_ccff_tail));

	grid_io_bottom grid_io_bottom_22__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[352:359]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_21__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[360:367]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_20__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[368:375]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_19__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[376:383]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_bottom grid_io_bottom_18__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[384:391]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_4_ccff_tail));

	grid_io_bottom grid_io_bottom_17__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[392:399]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_5_ccff_tail));

	grid_io_bottom grid_io_bottom_16__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[400:407]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_6_ccff_tail));

	grid_io_bottom grid_io_bottom_15__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[408:415]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_7_ccff_tail));

	grid_io_bottom grid_io_bottom_14__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[416:423]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_8_ccff_tail));

	grid_io_bottom grid_io_bottom_13__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[424:431]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_9_ccff_tail));

	grid_io_bottom grid_io_bottom_12__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[432:439]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_10_ccff_tail));

	grid_io_bottom grid_io_bottom_11__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[440:447]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_11_ccff_tail));

	grid_io_bottom grid_io_bottom_10__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[448:455]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_12_ccff_tail));

	grid_io_bottom grid_io_bottom_9__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[456:463]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_13_ccff_tail));

	grid_io_bottom grid_io_bottom_8__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[464:471]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_14_ccff_tail));

	grid_io_bottom grid_io_bottom_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[472:479]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_15_ccff_tail));

	grid_io_bottom grid_io_bottom_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[480:487]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_16_ccff_tail));

	grid_io_bottom grid_io_bottom_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[488:495]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_17_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[496:503]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_18_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[504:511]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_19_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[512:519]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_20_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[520:527]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_21_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[528:535]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[536:543]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[544:551]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[552:559]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[560:567]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__5__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[568:575]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_io_left grid_io_left_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[576:583]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_6_ccff_tail));

	grid_io_left grid_io_left_0__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[584:591]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_7_ccff_tail));

	grid_io_left grid_io_left_0__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[592:599]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_8_ccff_tail));

	grid_io_left grid_io_left_0__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[600:607]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__8_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_9_ccff_tail));

	grid_io_left grid_io_left_0__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[608:615]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__9_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_10_ccff_tail));

	grid_io_left grid_io_left_0__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[616:623]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__10_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_11_ccff_tail));

	grid_io_left grid_io_left_0__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[624:631]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__11_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_12_ccff_tail));

	grid_io_left grid_io_left_0__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[632:639]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__12_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_13_ccff_tail));

	grid_io_left grid_io_left_0__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[640:647]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__13_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_14_ccff_tail));

	grid_io_left grid_io_left_0__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[648:655]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__14_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_15_ccff_tail));

	grid_io_left grid_io_left_0__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[656:663]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__15_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_16_ccff_tail));

	grid_io_left grid_io_left_0__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[664:671]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__16_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_17_ccff_tail));

	grid_io_left grid_io_left_0__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[672:679]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__17_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_18_ccff_tail));

	grid_io_left grid_io_left_0__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[680:687]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__18_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_19_ccff_tail));

	grid_io_left grid_io_left_0__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[688:695]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__19_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_20_ccff_tail));

	grid_io_left grid_io_left_0__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[696:703]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__20_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_21_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_9__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_10__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_11__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_11__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_12__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_12__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_13__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_13__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_14__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_14__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_15__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_15__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_16__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_16__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_17__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_17__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_18__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_18__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_19__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_19__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_20__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_20__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_21__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_21__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__5__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_22__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_22__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_22__5__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_12_),
		.top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_7_),
		.left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_11_),
		.left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_15_),
		.left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_router grid_router_3__3_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_3__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_3__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_3__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_3__9_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_3__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_6__3_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_6__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_6__9_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_9__3_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_9__3__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_9__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_9__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	grid_router grid_router_9__9_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_9__9__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_1_));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:228]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:228]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_7_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__1_ sb_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_8_ccff_tail),
		.chany_top_out(sb_0__1__4_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__4_ccff_tail));

	sb_0__1_ sb_0__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_9_ccff_tail),
		.chany_top_out(sb_0__1__5_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__5_ccff_tail));

	sb_0__1_ sb_0__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__8_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_10_ccff_tail),
		.chany_top_out(sb_0__1__6_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__6_ccff_tail));

	sb_0__1_ sb_0__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__9_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_11_ccff_tail),
		.chany_top_out(sb_0__1__7_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__7_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__7_ccff_tail));

	sb_0__1_ sb_0__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__10_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_12_ccff_tail),
		.chany_top_out(sb_0__1__8_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__8_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__8_ccff_tail));

	sb_0__1_ sb_0__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__11_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__10_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_13_ccff_tail),
		.chany_top_out(sb_0__1__9_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__9_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__9_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__9_ccff_tail));

	sb_0__1_ sb_0__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__12_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__11_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_14_ccff_tail),
		.chany_top_out(sb_0__1__10_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__10_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__10_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__10_ccff_tail));

	sb_0__1_ sb_0__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__13_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__12_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_15_ccff_tail),
		.chany_top_out(sb_0__1__11_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__11_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__11_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__11_ccff_tail));

	sb_0__1_ sb_0__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__14_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__13_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_16_ccff_tail),
		.chany_top_out(sb_0__1__12_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__12_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__12_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__12_ccff_tail));

	sb_0__1_ sb_0__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__15_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__14_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_17_ccff_tail),
		.chany_top_out(sb_0__1__13_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__13_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__13_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__13_ccff_tail));

	sb_0__1_ sb_0__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__16_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__15_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_18_ccff_tail),
		.chany_top_out(sb_0__1__14_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__14_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__14_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__14_ccff_tail));

	sb_0__1_ sb_0__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__17_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__16_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_19_ccff_tail),
		.chany_top_out(sb_0__1__15_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__15_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__15_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__15_ccff_tail));

	sb_0__1_ sb_0__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__18_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__17_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_20_ccff_tail),
		.chany_top_out(sb_0__1__16_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__16_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__16_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__16_ccff_tail));

	sb_0__1_ sb_0__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__19_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__18_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_21_ccff_tail),
		.chany_top_out(sb_0__1__17_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__17_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__17_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__17_ccff_tail));

	sb_0__1_ sb_0__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__20_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:228]),
		.chany_bottom_in(cby_0__1__19_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_20_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__22__0_ccff_tail),
		.chany_top_out(sb_0__1__18_chany_top_out[0:228]),
		.chanx_right_out(sb_0__1__18_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__1__18_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__1__18_ccff_tail));

	sb_0__4_ sb_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__5__0_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__0_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_0__4__0_chany_top_out[0:228]),
		.chanx_right_out(sb_0__4__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__4__0_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__4__0_ccff_tail));

	sb_0__5_ sb_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__5__0_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_0__5__0_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_6_ccff_tail),
		.chany_top_out(sb_0__5__0_chany_top_out[0:228]),
		.chanx_right_out(sb_0__5__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__5__0_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__5__0_ccff_tail));

	sb_0__22_ sb_0__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__0_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__20_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_21_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__22__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_0__22__0_chany_bottom_out[0:228]),
		.ccff_tail(sb_0__22__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_21_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__21_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_20_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__39_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__57_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__78_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__0_ sb_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__96_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_top_out(sb_1__0__5_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__5_ccff_tail));

	sb_1__0_ sb_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__114_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.chany_top_out(sb_1__0__6_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__6_ccff_tail));

	sb_1__0_ sb_8__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__135_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__8_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__6_ccff_tail),
		.chany_top_out(sb_1__0__7_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__7_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__7_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__7_ccff_tail));

	sb_1__0_ sb_9__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__153_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__9_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__8_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__7_ccff_tail),
		.chany_top_out(sb_1__0__8_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__8_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__8_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__8_ccff_tail));

	sb_1__0_ sb_10__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__171_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__10_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__9_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__8_ccff_tail),
		.chany_top_out(sb_1__0__9_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__9_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__9_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__9_ccff_tail));

	sb_1__0_ sb_11__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__192_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__11_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__10_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__9_ccff_tail),
		.chany_top_out(sb_1__0__10_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__10_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__10_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__10_ccff_tail));

	sb_1__0_ sb_12__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__213_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__12_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__11_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__10_ccff_tail),
		.chany_top_out(sb_1__0__11_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__11_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__11_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__11_ccff_tail));

	sb_1__0_ sb_13__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__234_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__13_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__12_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__11_ccff_tail),
		.chany_top_out(sb_1__0__12_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__12_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__12_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__12_ccff_tail));

	sb_1__0_ sb_14__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__255_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__14_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__13_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__12_ccff_tail),
		.chany_top_out(sb_1__0__13_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__13_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__13_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__13_ccff_tail));

	sb_1__0_ sb_15__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__276_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__15_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__14_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__13_ccff_tail),
		.chany_top_out(sb_1__0__14_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__14_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__14_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__14_ccff_tail));

	sb_1__0_ sb_16__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__297_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__16_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__15_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__14_ccff_tail),
		.chany_top_out(sb_1__0__15_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__15_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__15_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__15_ccff_tail));

	sb_1__0_ sb_17__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__318_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__17_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__16_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__15_ccff_tail),
		.chany_top_out(sb_1__0__16_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__16_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__16_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__16_ccff_tail));

	sb_1__0_ sb_18__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__339_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__18_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__17_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__16_ccff_tail),
		.chany_top_out(sb_1__0__17_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__17_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__17_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__17_ccff_tail));

	sb_1__0_ sb_19__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__360_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__19_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__18_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__17_ccff_tail),
		.chany_top_out(sb_1__0__18_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__18_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__18_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__18_ccff_tail));

	sb_1__0_ sb_20__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__381_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__20_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__19_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__18_ccff_tail),
		.chany_top_out(sb_1__0__19_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__19_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__19_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__19_ccff_tail));

	sb_1__0_ sb_21__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__402_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__0__21_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__20_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__19_ccff_tail),
		.chany_top_out(sb_1__0__20_chany_top_out[0:228]),
		.chanx_right_out(sb_1__0__20_chanx_right_out[0:228]),
		.chanx_left_out(sb_1__0__20_chanx_left_out[0:228]),
		.ccff_tail(sb_1__0__20_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__19_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__20_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__21_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__0_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__22_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:228]),
		.ccff_head(cbx_1__5__0_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__23_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__20_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__24_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_1__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__25_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__2_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_1__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__26_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_1__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__27_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__22_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__1_ sb_1__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__28_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chany_top_out(sb_1__1__9_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__9_ccff_tail));

	sb_1__1_ sb_1__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__29_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__24_ccff_tail),
		.chany_top_out(sb_1__1__10_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__10_ccff_tail));

	sb_1__1_ sb_1__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__30_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__10_ccff_tail),
		.chany_top_out(sb_1__1__11_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__11_ccff_tail));

	sb_1__1_ sb_1__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__31_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__26_ccff_tail),
		.chany_top_out(sb_1__1__12_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__12_ccff_tail));

	sb_1__1_ sb_1__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__32_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__12_ccff_tail),
		.chany_top_out(sb_1__1__13_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__13_ccff_tail));

	sb_1__1_ sb_1__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__33_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__28_ccff_tail),
		.chany_top_out(sb_1__1__14_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__14_ccff_tail));

	sb_1__1_ sb_1__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__34_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__14_ccff_tail),
		.chany_top_out(sb_1__1__15_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__15_ccff_tail));

	sb_1__1_ sb_1__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__35_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__30_ccff_tail),
		.chany_top_out(sb_1__1__16_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__16_ccff_tail));

	sb_1__1_ sb_1__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__36_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__16_ccff_tail),
		.chany_top_out(sb_1__1__17_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__17_ccff_tail));

	sb_1__1_ sb_1__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__20_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__37_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__32_ccff_tail),
		.chany_top_out(sb_1__1__18_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:228]),
		.ccff_tail(ccff_tail));

	sb_1__1_ sb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__22_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__38_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__33_ccff_tail),
		.chany_top_out(sb_1__1__19_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__19_ccff_tail));

	sb_1__1_ sb_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__25_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__39_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__23_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__34_ccff_tail),
		.chany_top_out(sb_1__1__20_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__20_ccff_tail));

	sb_1__1_ sb_2__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__27_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__40_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__26_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chany_top_out(sb_1__1__21_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__21_ccff_tail));

	sb_1__1_ sb_2__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__28_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__41_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__27_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__36_ccff_tail),
		.chany_top_out(sb_1__1__22_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__22_ccff_tail));

	sb_1__1_ sb_2__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__29_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__42_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__28_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__9_ccff_tail),
		.chany_top_out(sb_1__1__23_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__23_ccff_tail));

	sb_1__1_ sb_2__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__30_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__43_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__29_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__38_ccff_tail),
		.chany_top_out(sb_1__1__24_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__24_ccff_tail));

	sb_1__1_ sb_2__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__31_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__44_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__30_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__11_ccff_tail),
		.chany_top_out(sb_1__1__25_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__25_ccff_tail));

	sb_1__1_ sb_2__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__32_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__45_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__31_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__40_ccff_tail),
		.chany_top_out(sb_1__1__26_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__26_ccff_tail));

	sb_1__1_ sb_2__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__33_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__46_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__32_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__13_ccff_tail),
		.chany_top_out(sb_1__1__27_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__27_ccff_tail));

	sb_1__1_ sb_2__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__34_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__47_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__33_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__42_ccff_tail),
		.chany_top_out(sb_1__1__28_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__28_ccff_tail));

	sb_1__1_ sb_2__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__35_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__48_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__34_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__15_ccff_tail),
		.chany_top_out(sb_1__1__29_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__29_ccff_tail));

	sb_1__1_ sb_2__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__36_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__49_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__35_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__44_ccff_tail),
		.chany_top_out(sb_1__1__30_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__30_ccff_tail));

	sb_1__1_ sb_2__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__37_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__50_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__36_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__17_ccff_tail),
		.chany_top_out(sb_1__1__31_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__31_ccff_tail));

	sb_1__1_ sb_2__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__38_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__51_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__37_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__46_ccff_tail),
		.chany_top_out(sb_1__1__32_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__32_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__40_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__52_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__38_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__47_ccff_tail),
		.chany_top_out(sb_1__1__33_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__33_ccff_tail));

	sb_1__1_ sb_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__43_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__56_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__39_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__51_ccff_tail),
		.chany_top_out(sb_1__1__34_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__34_ccff_tail));

	sb_1__1_ sb_3__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__45_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__59_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__40_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__21_ccff_tail),
		.chany_top_out(sb_1__1__35_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__35_ccff_tail));

	sb_1__1_ sb_3__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__46_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__60_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__41_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__55_ccff_tail),
		.chany_top_out(sb_1__1__36_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__36_ccff_tail));

	sb_1__1_ sb_3__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__47_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__61_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__42_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__23_ccff_tail),
		.chany_top_out(sb_1__1__37_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__37_ccff_tail));

	sb_1__1_ sb_3__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__48_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__62_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__43_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__57_ccff_tail),
		.chany_top_out(sb_1__1__38_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__38_ccff_tail));

	sb_1__1_ sb_3__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__49_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__63_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__44_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__25_ccff_tail),
		.chany_top_out(sb_1__1__39_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__39_ccff_tail));

	sb_1__1_ sb_3__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__50_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__64_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__45_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__59_ccff_tail),
		.chany_top_out(sb_1__1__40_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__40_ccff_tail));

	sb_1__1_ sb_3__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__51_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__65_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__46_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__27_ccff_tail),
		.chany_top_out(sb_1__1__41_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__41_ccff_tail));

	sb_1__1_ sb_3__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__52_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__66_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__47_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__61_ccff_tail),
		.chany_top_out(sb_1__1__42_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__42_ccff_tail));

	sb_1__1_ sb_3__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__53_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__67_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__48_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__29_ccff_tail),
		.chany_top_out(sb_1__1__43_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__43_ccff_tail));

	sb_1__1_ sb_3__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__54_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__68_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__49_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__63_ccff_tail),
		.chany_top_out(sb_1__1__44_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__44_ccff_tail));

	sb_1__1_ sb_3__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__55_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__69_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__50_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__31_ccff_tail),
		.chany_top_out(sb_1__1__45_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__45_ccff_tail));

	sb_1__1_ sb_3__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__56_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__70_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__51_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__65_ccff_tail),
		.chany_top_out(sb_1__1__46_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__46_ccff_tail));

	sb_1__1_ sb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__58_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__71_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__57_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__52_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__66_ccff_tail),
		.chany_top_out(sb_1__1__47_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__47_ccff_tail));

	sb_1__1_ sb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__59_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__72_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__58_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__53_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__0_ccff_tail),
		.chany_top_out(sb_1__1__48_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__48_ccff_tail));

	sb_1__1_ sb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__60_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__73_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__59_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__54_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__3_ccff_tail),
		.chany_top_out(sb_1__1__49_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__49_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__49_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__49_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__49_ccff_tail));

	sb_1__1_ sb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__62_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__74_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__61_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__55_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__1_ccff_tail),
		.chany_top_out(sb_1__1__50_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__50_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__50_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__50_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__50_ccff_tail));

	sb_1__1_ sb_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__63_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__75_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__62_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__56_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__67_ccff_tail),
		.chany_top_out(sb_1__1__51_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__51_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__51_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__51_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__51_ccff_tail));

	sb_1__1_ sb_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__64_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__76_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__63_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__57_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__2_ccff_tail),
		.chany_top_out(sb_1__1__52_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__52_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__52_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__52_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__52_ccff_tail));

	sb_1__1_ sb_4__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__65_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__77_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__64_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__58_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__5_ccff_tail),
		.chany_top_out(sb_1__1__53_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__53_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__53_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__53_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__53_ccff_tail));

	sb_1__1_ sb_4__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__66_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__78_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__65_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__59_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__35_ccff_tail),
		.chany_top_out(sb_1__1__54_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__54_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__54_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__54_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__54_ccff_tail));

	sb_1__1_ sb_4__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__67_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__79_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__66_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__60_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__69_ccff_tail),
		.chany_top_out(sb_1__1__55_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__55_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__55_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__55_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__55_ccff_tail));

	sb_1__1_ sb_4__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__68_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__80_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__67_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__61_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__37_ccff_tail),
		.chany_top_out(sb_1__1__56_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__56_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__56_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__56_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__56_ccff_tail));

	sb_1__1_ sb_4__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__69_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__81_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__68_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__62_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__71_ccff_tail),
		.chany_top_out(sb_1__1__57_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__57_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__57_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__57_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__57_ccff_tail));

	sb_1__1_ sb_4__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__70_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__82_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__69_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__63_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__39_ccff_tail),
		.chany_top_out(sb_1__1__58_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__58_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__58_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__58_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__58_ccff_tail));

	sb_1__1_ sb_4__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__71_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__83_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__70_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__64_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__73_ccff_tail),
		.chany_top_out(sb_1__1__59_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__59_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__59_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__59_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__59_ccff_tail));

	sb_1__1_ sb_4__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__72_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__84_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__71_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__65_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__41_ccff_tail),
		.chany_top_out(sb_1__1__60_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__60_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__60_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__60_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__60_ccff_tail));

	sb_1__1_ sb_4__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__73_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__85_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__72_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__66_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__75_ccff_tail),
		.chany_top_out(sb_1__1__61_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__61_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__61_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__61_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__61_ccff_tail));

	sb_1__1_ sb_4__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__74_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__86_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__73_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__67_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__43_ccff_tail),
		.chany_top_out(sb_1__1__62_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__62_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__62_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__62_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__62_ccff_tail));

	sb_1__1_ sb_4__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__75_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__87_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__74_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__68_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__77_ccff_tail),
		.chany_top_out(sb_1__1__63_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__63_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__63_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__63_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__63_ccff_tail));

	sb_1__1_ sb_4__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__76_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__88_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__75_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__69_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__45_ccff_tail),
		.chany_top_out(sb_1__1__64_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__64_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__64_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__64_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__64_ccff_tail));

	sb_1__1_ sb_4__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__77_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__89_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__76_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__70_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__79_ccff_tail),
		.chany_top_out(sb_1__1__65_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__65_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__65_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__65_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__65_ccff_tail));

	sb_1__1_ sb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__79_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__90_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__78_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__71_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__80_ccff_tail),
		.chany_top_out(sb_1__1__66_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__66_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__66_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__66_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__66_ccff_tail));

	sb_1__1_ sb_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__82_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__91_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__81_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__75_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__81_ccff_tail),
		.chany_top_out(sb_1__1__67_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__67_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__67_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__67_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__67_ccff_tail));

	sb_1__1_ sb_5__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__84_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__92_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__83_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__78_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__54_ccff_tail),
		.chany_top_out(sb_1__1__68_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__68_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__68_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__68_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__68_ccff_tail));

	sb_1__1_ sb_5__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__85_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__93_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__84_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__79_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__83_ccff_tail),
		.chany_top_out(sb_1__1__69_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__69_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__69_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__69_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__69_ccff_tail));

	sb_1__1_ sb_5__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__86_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__94_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__85_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__80_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__56_ccff_tail),
		.chany_top_out(sb_1__1__70_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__70_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__70_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__70_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__70_ccff_tail));

	sb_1__1_ sb_5__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__87_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__95_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__86_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__81_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__85_ccff_tail),
		.chany_top_out(sb_1__1__71_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__71_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__71_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__71_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__71_ccff_tail));

	sb_1__1_ sb_5__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__88_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__96_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__87_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__82_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__58_ccff_tail),
		.chany_top_out(sb_1__1__72_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__72_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__72_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__72_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__72_ccff_tail));

	sb_1__1_ sb_5__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__89_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__97_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__88_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__83_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__87_ccff_tail),
		.chany_top_out(sb_1__1__73_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__73_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__73_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__73_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__73_ccff_tail));

	sb_1__1_ sb_5__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__90_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__98_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__89_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__84_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__60_ccff_tail),
		.chany_top_out(sb_1__1__74_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__74_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__74_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__74_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__74_ccff_tail));

	sb_1__1_ sb_5__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__91_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__99_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__90_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__85_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__89_ccff_tail),
		.chany_top_out(sb_1__1__75_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__75_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__75_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__75_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__75_ccff_tail));

	sb_1__1_ sb_5__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__92_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__100_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__91_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__86_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__62_ccff_tail),
		.chany_top_out(sb_1__1__76_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__76_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__76_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__76_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__76_ccff_tail));

	sb_1__1_ sb_5__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__93_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__101_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__92_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__87_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__91_ccff_tail),
		.chany_top_out(sb_1__1__77_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__77_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__77_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__77_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__77_ccff_tail));

	sb_1__1_ sb_5__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__94_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__102_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__93_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__88_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__64_ccff_tail),
		.chany_top_out(sb_1__1__78_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__78_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__78_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__78_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__78_ccff_tail));

	sb_1__1_ sb_5__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__95_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__103_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__94_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__89_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__93_ccff_tail),
		.chany_top_out(sb_1__1__79_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__79_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__79_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__79_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__79_ccff_tail));

	sb_1__1_ sb_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__97_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__104_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__96_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__90_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__94_ccff_tail),
		.chany_top_out(sb_1__1__80_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__80_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__80_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__80_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__80_ccff_tail));

	sb_1__1_ sb_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__100_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__108_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__99_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__91_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__98_ccff_tail),
		.chany_top_out(sb_1__1__81_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__81_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__81_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__81_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__81_ccff_tail));

	sb_1__1_ sb_6__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__102_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__111_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__101_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__92_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__68_ccff_tail),
		.chany_top_out(sb_1__1__82_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__82_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__82_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__82_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__82_ccff_tail));

	sb_1__1_ sb_6__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__103_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__112_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__102_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__93_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__102_ccff_tail),
		.chany_top_out(sb_1__1__83_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__83_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__83_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__83_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__83_ccff_tail));

	sb_1__1_ sb_6__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__104_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__113_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__103_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__94_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__70_ccff_tail),
		.chany_top_out(sb_1__1__84_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__84_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__84_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__84_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__84_ccff_tail));

	sb_1__1_ sb_6__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__105_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__114_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__104_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__95_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__104_ccff_tail),
		.chany_top_out(sb_1__1__85_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__85_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__85_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__85_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__85_ccff_tail));

	sb_1__1_ sb_6__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__106_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__115_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__105_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__96_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__72_ccff_tail),
		.chany_top_out(sb_1__1__86_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__86_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__86_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__86_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__86_ccff_tail));

	sb_1__1_ sb_6__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__107_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__116_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__106_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__97_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__106_ccff_tail),
		.chany_top_out(sb_1__1__87_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__87_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__87_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__87_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__87_ccff_tail));

	sb_1__1_ sb_6__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__108_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__117_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__107_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__98_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__74_ccff_tail),
		.chany_top_out(sb_1__1__88_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__88_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__88_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__88_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__88_ccff_tail));

	sb_1__1_ sb_6__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__109_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__118_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__108_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__99_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__108_ccff_tail),
		.chany_top_out(sb_1__1__89_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__89_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__89_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__89_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__89_ccff_tail));

	sb_1__1_ sb_6__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__110_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__119_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__109_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__100_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__76_ccff_tail),
		.chany_top_out(sb_1__1__90_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__90_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__90_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__90_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__90_ccff_tail));

	sb_1__1_ sb_6__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__111_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__120_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__110_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__101_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__110_ccff_tail),
		.chany_top_out(sb_1__1__91_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__91_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__91_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__91_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__91_ccff_tail));

	sb_1__1_ sb_6__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__112_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__121_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__111_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__102_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__78_ccff_tail),
		.chany_top_out(sb_1__1__92_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__92_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__92_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__92_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__92_ccff_tail));

	sb_1__1_ sb_6__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__113_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__122_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__112_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__103_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__112_ccff_tail),
		.chany_top_out(sb_1__1__93_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__93_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__93_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__93_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__93_ccff_tail));

	sb_1__1_ sb_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__115_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__123_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__114_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__104_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__113_ccff_tail),
		.chany_top_out(sb_1__1__94_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__94_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__94_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__94_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__94_ccff_tail));

	sb_1__1_ sb_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__116_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__124_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__115_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__105_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__3_ccff_tail),
		.chany_top_out(sb_1__1__95_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__95_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__95_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__95_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__95_ccff_tail));

	sb_1__1_ sb_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__117_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__125_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__116_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__106_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__6_ccff_tail),
		.chany_top_out(sb_1__1__96_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__96_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__96_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__96_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__96_ccff_tail));

	sb_1__1_ sb_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__119_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__126_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__118_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__107_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__4_ccff_tail),
		.chany_top_out(sb_1__1__97_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__97_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__97_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__97_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__97_ccff_tail));

	sb_1__1_ sb_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__120_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__127_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__119_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__108_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__114_ccff_tail),
		.chany_top_out(sb_1__1__98_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__98_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__98_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__98_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__98_ccff_tail));

	sb_1__1_ sb_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__121_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__128_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__120_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__109_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__5_ccff_tail),
		.chany_top_out(sb_1__1__99_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__99_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__99_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__99_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__99_ccff_tail));

	sb_1__1_ sb_7__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__122_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__129_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__121_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__110_chanx_right_out[0:228]),
		.ccff_head(sb_2__3__8_ccff_tail),
		.chany_top_out(sb_1__1__100_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__100_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__100_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__100_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__100_ccff_tail));

	sb_1__1_ sb_7__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__123_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__130_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__122_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__111_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__82_ccff_tail),
		.chany_top_out(sb_1__1__101_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__101_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__101_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__101_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__101_ccff_tail));

	sb_1__1_ sb_7__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__124_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__131_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__123_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__112_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__116_ccff_tail),
		.chany_top_out(sb_1__1__102_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__102_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__102_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__102_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__102_ccff_tail));

	sb_1__1_ sb_7__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__125_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__132_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__124_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__113_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__84_ccff_tail),
		.chany_top_out(sb_1__1__103_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__103_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__103_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__103_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__103_ccff_tail));

	sb_1__1_ sb_7__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__126_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__133_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__125_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__114_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__118_ccff_tail),
		.chany_top_out(sb_1__1__104_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__104_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__104_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__104_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__104_ccff_tail));

	sb_1__1_ sb_7__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__127_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__134_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__126_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__115_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__86_ccff_tail),
		.chany_top_out(sb_1__1__105_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__105_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__105_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__105_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__105_ccff_tail));

	sb_1__1_ sb_7__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__128_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__135_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__127_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__116_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__120_ccff_tail),
		.chany_top_out(sb_1__1__106_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__106_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__106_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__106_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__106_ccff_tail));

	sb_1__1_ sb_7__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__129_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__136_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__128_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__117_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__88_ccff_tail),
		.chany_top_out(sb_1__1__107_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__107_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__107_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__107_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__107_ccff_tail));

	sb_1__1_ sb_7__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__130_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__137_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__129_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__118_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__122_ccff_tail),
		.chany_top_out(sb_1__1__108_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__108_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__108_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__108_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__108_ccff_tail));

	sb_1__1_ sb_7__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__131_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__138_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__130_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__119_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__90_ccff_tail),
		.chany_top_out(sb_1__1__109_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__109_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__109_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__109_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__109_ccff_tail));

	sb_1__1_ sb_7__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__132_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__139_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__131_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__120_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__124_ccff_tail),
		.chany_top_out(sb_1__1__110_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__110_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__110_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__110_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__110_ccff_tail));

	sb_1__1_ sb_7__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__133_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__140_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__132_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__121_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__92_ccff_tail),
		.chany_top_out(sb_1__1__111_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__111_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__111_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__111_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__111_ccff_tail));

	sb_1__1_ sb_7__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__134_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__141_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__133_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__122_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__126_ccff_tail),
		.chany_top_out(sb_1__1__112_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__112_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__112_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__112_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__112_ccff_tail));

	sb_1__1_ sb_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__136_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__142_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__135_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__123_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__127_ccff_tail),
		.chany_top_out(sb_1__1__113_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__113_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__113_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__113_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__113_ccff_tail));

	sb_1__1_ sb_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__139_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__143_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__138_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__127_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__128_ccff_tail),
		.chany_top_out(sb_1__1__114_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__114_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__114_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__114_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__114_ccff_tail));

	sb_1__1_ sb_8__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__141_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__144_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__140_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__130_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__101_ccff_tail),
		.chany_top_out(sb_1__1__115_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__115_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__115_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__115_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__115_ccff_tail));

	sb_1__1_ sb_8__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__142_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__145_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__141_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__131_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__130_ccff_tail),
		.chany_top_out(sb_1__1__116_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__116_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__116_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__116_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__116_ccff_tail));

	sb_1__1_ sb_8__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__143_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__146_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__142_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__132_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__103_ccff_tail),
		.chany_top_out(sb_1__1__117_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__117_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__117_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__117_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__117_ccff_tail));

	sb_1__1_ sb_8__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__144_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__147_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__143_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__133_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__132_ccff_tail),
		.chany_top_out(sb_1__1__118_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__118_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__118_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__118_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__118_ccff_tail));

	sb_1__1_ sb_8__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__145_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__148_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__144_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__134_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__105_ccff_tail),
		.chany_top_out(sb_1__1__119_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__119_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__119_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__119_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__119_ccff_tail));

	sb_1__1_ sb_8__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__146_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__149_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__145_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__135_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__134_ccff_tail),
		.chany_top_out(sb_1__1__120_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__120_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__120_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__120_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__120_ccff_tail));

	sb_1__1_ sb_8__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__147_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__150_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__146_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__136_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__107_ccff_tail),
		.chany_top_out(sb_1__1__121_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__121_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__121_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__121_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__121_ccff_tail));

	sb_1__1_ sb_8__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__148_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__151_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__147_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__137_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__136_ccff_tail),
		.chany_top_out(sb_1__1__122_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__122_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__122_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__122_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__122_ccff_tail));

	sb_1__1_ sb_8__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__149_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__152_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__148_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__138_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__109_ccff_tail),
		.chany_top_out(sb_1__1__123_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__123_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__123_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__123_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__123_ccff_tail));

	sb_1__1_ sb_8__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__150_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__153_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__149_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__139_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__138_ccff_tail),
		.chany_top_out(sb_1__1__124_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__124_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__124_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__124_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__124_ccff_tail));

	sb_1__1_ sb_8__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__151_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__154_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__150_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__140_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__111_ccff_tail),
		.chany_top_out(sb_1__1__125_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__125_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__125_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__125_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__125_ccff_tail));

	sb_1__1_ sb_8__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__152_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__155_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__151_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__141_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__140_ccff_tail),
		.chany_top_out(sb_1__1__126_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__126_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__126_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__126_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__126_ccff_tail));

	sb_1__1_ sb_9__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__154_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__156_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__153_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__142_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__141_ccff_tail),
		.chany_top_out(sb_1__1__127_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__127_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__127_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__127_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__127_ccff_tail));

	sb_1__1_ sb_9__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__157_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__160_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__156_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__143_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__145_ccff_tail),
		.chany_top_out(sb_1__1__128_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__128_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__128_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__128_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__128_ccff_tail));

	sb_1__1_ sb_9__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__159_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__163_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__158_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__144_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__115_ccff_tail),
		.chany_top_out(sb_1__1__129_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__129_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__129_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__129_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__129_ccff_tail));

	sb_1__1_ sb_9__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__160_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__164_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__159_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__145_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__149_ccff_tail),
		.chany_top_out(sb_1__1__130_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__130_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__130_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__130_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__130_ccff_tail));

	sb_1__1_ sb_9__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__161_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__165_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__160_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__146_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__117_ccff_tail),
		.chany_top_out(sb_1__1__131_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__131_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__131_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__131_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__131_ccff_tail));

	sb_1__1_ sb_9__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__162_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__166_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__161_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__147_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__151_ccff_tail),
		.chany_top_out(sb_1__1__132_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__132_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__132_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__132_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__132_ccff_tail));

	sb_1__1_ sb_9__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__163_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__167_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__162_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__148_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__119_ccff_tail),
		.chany_top_out(sb_1__1__133_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__133_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__133_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__133_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__133_ccff_tail));

	sb_1__1_ sb_9__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__164_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__168_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__163_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__149_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__153_ccff_tail),
		.chany_top_out(sb_1__1__134_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__134_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__134_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__134_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__134_ccff_tail));

	sb_1__1_ sb_9__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__165_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__169_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__164_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__150_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__121_ccff_tail),
		.chany_top_out(sb_1__1__135_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__135_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__135_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__135_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__135_ccff_tail));

	sb_1__1_ sb_9__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__166_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__170_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__165_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__151_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__155_ccff_tail),
		.chany_top_out(sb_1__1__136_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__136_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__136_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__136_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__136_ccff_tail));

	sb_1__1_ sb_9__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__167_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__171_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__166_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__152_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__123_ccff_tail),
		.chany_top_out(sb_1__1__137_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__137_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__137_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__137_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__137_ccff_tail));

	sb_1__1_ sb_9__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__168_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__172_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__167_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__153_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__157_ccff_tail),
		.chany_top_out(sb_1__1__138_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__138_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__138_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__138_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__138_ccff_tail));

	sb_1__1_ sb_9__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__169_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__173_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__168_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__154_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__125_ccff_tail),
		.chany_top_out(sb_1__1__139_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__139_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__139_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__139_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__139_ccff_tail));

	sb_1__1_ sb_9__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__170_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__174_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__169_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__155_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__159_ccff_tail),
		.chany_top_out(sb_1__1__140_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__140_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__140_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__140_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__140_ccff_tail));

	sb_1__1_ sb_10__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__172_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__175_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__171_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__156_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__160_ccff_tail),
		.chany_top_out(sb_1__1__141_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__141_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__141_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__141_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__141_ccff_tail));

	sb_1__1_ sb_10__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__173_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__176_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__172_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__157_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__6_ccff_tail),
		.chany_top_out(sb_1__1__142_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__142_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__142_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__142_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__142_ccff_tail));

	sb_1__1_ sb_10__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__174_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__177_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__173_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__158_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__162_ccff_tail),
		.chany_top_out(sb_1__1__143_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__143_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__143_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__143_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__143_ccff_tail));

	sb_1__1_ sb_10__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__176_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__178_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__175_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__159_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__7_ccff_tail),
		.chany_top_out(sb_1__1__144_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__144_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__144_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__144_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__144_ccff_tail));

	sb_1__1_ sb_10__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__177_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__179_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__176_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__160_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__164_ccff_tail),
		.chany_top_out(sb_1__1__145_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__145_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__145_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__145_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__145_ccff_tail));

	sb_1__1_ sb_10__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__178_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__180_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__177_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__161_chanx_right_out[0:228]),
		.ccff_head(cby_3__3__8_ccff_tail),
		.chany_top_out(sb_1__1__146_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__146_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__146_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__146_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__146_ccff_tail));

	sb_1__1_ sb_10__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__179_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__181_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__178_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__162_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__166_ccff_tail),
		.chany_top_out(sb_1__1__147_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__147_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__147_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__147_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__147_ccff_tail));

	sb_1__1_ sb_10__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__180_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__182_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__179_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__163_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__129_ccff_tail),
		.chany_top_out(sb_1__1__148_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__148_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__148_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__148_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__148_ccff_tail));

	sb_1__1_ sb_10__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__181_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__183_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__180_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__164_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__168_ccff_tail),
		.chany_top_out(sb_1__1__149_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__149_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__149_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__149_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__149_ccff_tail));

	sb_1__1_ sb_10__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__182_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__184_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__181_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__165_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__131_ccff_tail),
		.chany_top_out(sb_1__1__150_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__150_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__150_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__150_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__150_ccff_tail));

	sb_1__1_ sb_10__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__183_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__185_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__182_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__166_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__170_ccff_tail),
		.chany_top_out(sb_1__1__151_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__151_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__151_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__151_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__151_ccff_tail));

	sb_1__1_ sb_10__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__184_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__186_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__183_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__167_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__133_ccff_tail),
		.chany_top_out(sb_1__1__152_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__152_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__152_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__152_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__152_ccff_tail));

	sb_1__1_ sb_10__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__185_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__187_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__184_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__168_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__172_ccff_tail),
		.chany_top_out(sb_1__1__153_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__153_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__153_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__153_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__153_ccff_tail));

	sb_1__1_ sb_10__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__186_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__188_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__185_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__169_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__135_ccff_tail),
		.chany_top_out(sb_1__1__154_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__154_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__154_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__154_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__154_ccff_tail));

	sb_1__1_ sb_10__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__187_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__189_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__186_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__170_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__174_ccff_tail),
		.chany_top_out(sb_1__1__155_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__155_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__155_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__155_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__155_ccff_tail));

	sb_1__1_ sb_10__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__188_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__190_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__187_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__171_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__137_ccff_tail),
		.chany_top_out(sb_1__1__156_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__156_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__156_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__156_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__156_ccff_tail));

	sb_1__1_ sb_10__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__189_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__191_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__188_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__172_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__176_ccff_tail),
		.chany_top_out(sb_1__1__157_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__157_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__157_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__157_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__157_ccff_tail));

	sb_1__1_ sb_10__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__190_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__192_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__189_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__173_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__139_ccff_tail),
		.chany_top_out(sb_1__1__158_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__158_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__158_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__158_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__158_ccff_tail));

	sb_1__1_ sb_10__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__191_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__193_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__190_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__174_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__178_ccff_tail),
		.chany_top_out(sb_1__1__159_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__159_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__159_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__159_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__159_ccff_tail));

	sb_1__1_ sb_11__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__193_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__194_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__192_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__175_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__179_ccff_tail),
		.chany_top_out(sb_1__1__160_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__160_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__160_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__160_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__160_ccff_tail));

	sb_1__1_ sb_11__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__194_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__195_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__193_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__176_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__142_ccff_tail),
		.chany_top_out(sb_1__1__161_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__161_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__161_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__161_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__161_ccff_tail));

	sb_1__1_ sb_11__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__195_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__196_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__194_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__177_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__181_ccff_tail),
		.chany_top_out(sb_1__1__162_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__162_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__162_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__162_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__162_ccff_tail));

	sb_1__1_ sb_11__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__197_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__197_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__196_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__178_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__144_ccff_tail),
		.chany_top_out(sb_1__1__163_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__163_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__163_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__163_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__163_ccff_tail));

	sb_1__1_ sb_11__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__198_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__198_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__197_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__179_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__183_ccff_tail),
		.chany_top_out(sb_1__1__164_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__164_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__164_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__164_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__164_ccff_tail));

	sb_1__1_ sb_11__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__199_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__199_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__198_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__180_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__146_ccff_tail),
		.chany_top_out(sb_1__1__165_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__165_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__165_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__165_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__165_ccff_tail));

	sb_1__1_ sb_11__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__200_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__200_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__199_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__181_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__185_ccff_tail),
		.chany_top_out(sb_1__1__166_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__166_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__166_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__166_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__166_ccff_tail));

	sb_1__1_ sb_11__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__201_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__201_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__200_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__182_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__148_ccff_tail),
		.chany_top_out(sb_1__1__167_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__167_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__167_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__167_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__167_ccff_tail));

	sb_1__1_ sb_11__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__202_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__202_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__201_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__183_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__187_ccff_tail),
		.chany_top_out(sb_1__1__168_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__168_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__168_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__168_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__168_ccff_tail));

	sb_1__1_ sb_11__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__203_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__203_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__202_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__184_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__150_ccff_tail),
		.chany_top_out(sb_1__1__169_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__169_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__169_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__169_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__169_ccff_tail));

	sb_1__1_ sb_11__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__204_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__204_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__203_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__185_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__189_ccff_tail),
		.chany_top_out(sb_1__1__170_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__170_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__170_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__170_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__170_ccff_tail));

	sb_1__1_ sb_11__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__205_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__205_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__204_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__186_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__152_ccff_tail),
		.chany_top_out(sb_1__1__171_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__171_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__171_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__171_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__171_ccff_tail));

	sb_1__1_ sb_11__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__206_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__206_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__205_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__187_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__191_ccff_tail),
		.chany_top_out(sb_1__1__172_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__172_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__172_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__172_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__172_ccff_tail));

	sb_1__1_ sb_11__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__207_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__207_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__206_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__188_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__154_ccff_tail),
		.chany_top_out(sb_1__1__173_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__173_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__173_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__173_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__173_ccff_tail));

	sb_1__1_ sb_11__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__208_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__208_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__207_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__189_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__193_ccff_tail),
		.chany_top_out(sb_1__1__174_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__174_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__174_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__174_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__174_ccff_tail));

	sb_1__1_ sb_11__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__209_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__209_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__208_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__190_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__156_ccff_tail),
		.chany_top_out(sb_1__1__175_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__175_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__175_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__175_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__175_ccff_tail));

	sb_1__1_ sb_11__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__210_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__210_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__209_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__191_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__195_ccff_tail),
		.chany_top_out(sb_1__1__176_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__176_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__176_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__176_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__176_ccff_tail));

	sb_1__1_ sb_11__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__211_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__211_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__210_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__192_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__158_ccff_tail),
		.chany_top_out(sb_1__1__177_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__177_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__177_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__177_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__177_ccff_tail));

	sb_1__1_ sb_11__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__212_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__212_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__211_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__193_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__197_ccff_tail),
		.chany_top_out(sb_1__1__178_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__178_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__178_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__178_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__178_ccff_tail));

	sb_1__1_ sb_12__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__214_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__213_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__213_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__194_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__198_ccff_tail),
		.chany_top_out(sb_1__1__179_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__179_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__179_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__179_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__179_ccff_tail));

	sb_1__1_ sb_12__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__215_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__214_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__214_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__195_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__161_ccff_tail),
		.chany_top_out(sb_1__1__180_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__180_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__180_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__180_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__180_ccff_tail));

	sb_1__1_ sb_12__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__216_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__215_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__215_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__196_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__200_ccff_tail),
		.chany_top_out(sb_1__1__181_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__181_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__181_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__181_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__181_ccff_tail));

	sb_1__1_ sb_12__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__218_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__216_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__217_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__197_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__163_ccff_tail),
		.chany_top_out(sb_1__1__182_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__182_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__182_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__182_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__182_ccff_tail));

	sb_1__1_ sb_12__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__219_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__217_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__218_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__198_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__202_ccff_tail),
		.chany_top_out(sb_1__1__183_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__183_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__183_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__183_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__183_ccff_tail));

	sb_1__1_ sb_12__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__220_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__218_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__219_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__199_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__165_ccff_tail),
		.chany_top_out(sb_1__1__184_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__184_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__184_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__184_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__184_ccff_tail));

	sb_1__1_ sb_12__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__221_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__219_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__220_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__200_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__204_ccff_tail),
		.chany_top_out(sb_1__1__185_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__185_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__185_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__185_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__185_ccff_tail));

	sb_1__1_ sb_12__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__222_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__220_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__221_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__201_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__167_ccff_tail),
		.chany_top_out(sb_1__1__186_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__186_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__186_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__186_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__186_ccff_tail));

	sb_1__1_ sb_12__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__223_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__221_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__222_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__202_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__206_ccff_tail),
		.chany_top_out(sb_1__1__187_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__187_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__187_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__187_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__187_ccff_tail));

	sb_1__1_ sb_12__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__224_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__222_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__223_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__203_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__169_ccff_tail),
		.chany_top_out(sb_1__1__188_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__188_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__188_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__188_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__188_ccff_tail));

	sb_1__1_ sb_12__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__225_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__223_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__224_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__204_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__208_ccff_tail),
		.chany_top_out(sb_1__1__189_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__189_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__189_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__189_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__189_ccff_tail));

	sb_1__1_ sb_12__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__226_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__224_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__225_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__205_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__171_ccff_tail),
		.chany_top_out(sb_1__1__190_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__190_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__190_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__190_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__190_ccff_tail));

	sb_1__1_ sb_12__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__227_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__225_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__226_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__206_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__210_ccff_tail),
		.chany_top_out(sb_1__1__191_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__191_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__191_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__191_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__191_ccff_tail));

	sb_1__1_ sb_12__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__228_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__226_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__227_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__207_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__173_ccff_tail),
		.chany_top_out(sb_1__1__192_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__192_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__192_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__192_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__192_ccff_tail));

	sb_1__1_ sb_12__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__229_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__227_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__228_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__208_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__212_ccff_tail),
		.chany_top_out(sb_1__1__193_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__193_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__193_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__193_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__193_ccff_tail));

	sb_1__1_ sb_12__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__230_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__228_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__229_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__209_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__175_ccff_tail),
		.chany_top_out(sb_1__1__194_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__194_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__194_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__194_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__194_ccff_tail));

	sb_1__1_ sb_12__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__231_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__229_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__230_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__210_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__214_ccff_tail),
		.chany_top_out(sb_1__1__195_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__195_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__195_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__195_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__195_ccff_tail));

	sb_1__1_ sb_12__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__232_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__230_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__231_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__211_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__177_ccff_tail),
		.chany_top_out(sb_1__1__196_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__196_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__196_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__196_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__196_ccff_tail));

	sb_1__1_ sb_12__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__233_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__231_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__232_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__212_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__216_ccff_tail),
		.chany_top_out(sb_1__1__197_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__197_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__197_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__197_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__197_ccff_tail));

	sb_1__1_ sb_13__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__235_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__232_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__234_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__213_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__217_ccff_tail),
		.chany_top_out(sb_1__1__198_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__198_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__198_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__198_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__198_ccff_tail));

	sb_1__1_ sb_13__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__236_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__233_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__235_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__214_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__180_ccff_tail),
		.chany_top_out(sb_1__1__199_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__199_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__199_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__199_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__199_ccff_tail));

	sb_1__1_ sb_13__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__237_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__234_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__236_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__215_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__219_ccff_tail),
		.chany_top_out(sb_1__1__200_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__200_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__200_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__200_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__200_ccff_tail));

	sb_1__1_ sb_13__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__239_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__235_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__238_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__216_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__182_ccff_tail),
		.chany_top_out(sb_1__1__201_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__201_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__201_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__201_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__201_ccff_tail));

	sb_1__1_ sb_13__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__240_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__236_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__239_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__217_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__221_ccff_tail),
		.chany_top_out(sb_1__1__202_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__202_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__202_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__202_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__202_ccff_tail));

	sb_1__1_ sb_13__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__241_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__237_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__240_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__218_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__184_ccff_tail),
		.chany_top_out(sb_1__1__203_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__203_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__203_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__203_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__203_ccff_tail));

	sb_1__1_ sb_13__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__242_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__238_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__241_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__219_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__223_ccff_tail),
		.chany_top_out(sb_1__1__204_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__204_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__204_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__204_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__204_ccff_tail));

	sb_1__1_ sb_13__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__243_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__239_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__242_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__220_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__186_ccff_tail),
		.chany_top_out(sb_1__1__205_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__205_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__205_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__205_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__205_ccff_tail));

	sb_1__1_ sb_13__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__244_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__240_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__243_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__221_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__225_ccff_tail),
		.chany_top_out(sb_1__1__206_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__206_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__206_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__206_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__206_ccff_tail));

	sb_1__1_ sb_13__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__245_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__241_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__244_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__222_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__188_ccff_tail),
		.chany_top_out(sb_1__1__207_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__207_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__207_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__207_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__207_ccff_tail));

	sb_1__1_ sb_13__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__246_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__242_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__245_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__223_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__227_ccff_tail),
		.chany_top_out(sb_1__1__208_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__208_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__208_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__208_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__208_ccff_tail));

	sb_1__1_ sb_13__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__247_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__243_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__246_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__224_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__190_ccff_tail),
		.chany_top_out(sb_1__1__209_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__209_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__209_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__209_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__209_ccff_tail));

	sb_1__1_ sb_13__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__248_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__244_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__247_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__225_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__229_ccff_tail),
		.chany_top_out(sb_1__1__210_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__210_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__210_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__210_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__210_ccff_tail));

	sb_1__1_ sb_13__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__249_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__245_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__248_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__226_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__192_ccff_tail),
		.chany_top_out(sb_1__1__211_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__211_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__211_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__211_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__211_ccff_tail));

	sb_1__1_ sb_13__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__250_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__246_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__249_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__227_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__231_ccff_tail),
		.chany_top_out(sb_1__1__212_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__212_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__212_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__212_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__212_ccff_tail));

	sb_1__1_ sb_13__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__251_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__247_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__250_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__228_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__194_ccff_tail),
		.chany_top_out(sb_1__1__213_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__213_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__213_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__213_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__213_ccff_tail));

	sb_1__1_ sb_13__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__252_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__248_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__251_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__229_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__233_ccff_tail),
		.chany_top_out(sb_1__1__214_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__214_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__214_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__214_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__214_ccff_tail));

	sb_1__1_ sb_13__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__253_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__249_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__252_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__230_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__196_ccff_tail),
		.chany_top_out(sb_1__1__215_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__215_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__215_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__215_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__215_ccff_tail));

	sb_1__1_ sb_13__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__254_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__250_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__253_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__231_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__235_ccff_tail),
		.chany_top_out(sb_1__1__216_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__216_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__216_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__216_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__216_ccff_tail));

	sb_1__1_ sb_14__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__256_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__251_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__255_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__232_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__236_ccff_tail),
		.chany_top_out(sb_1__1__217_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__217_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__217_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__217_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__217_ccff_tail));

	sb_1__1_ sb_14__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__257_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__252_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__256_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__233_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__199_ccff_tail),
		.chany_top_out(sb_1__1__218_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__218_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__218_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__218_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__218_ccff_tail));

	sb_1__1_ sb_14__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__258_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__253_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__257_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__234_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__238_ccff_tail),
		.chany_top_out(sb_1__1__219_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__219_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__219_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__219_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__219_ccff_tail));

	sb_1__1_ sb_14__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__260_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__254_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__259_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__235_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__201_ccff_tail),
		.chany_top_out(sb_1__1__220_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__220_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__220_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__220_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__220_ccff_tail));

	sb_1__1_ sb_14__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__261_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__255_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__260_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__236_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__240_ccff_tail),
		.chany_top_out(sb_1__1__221_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__221_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__221_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__221_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__221_ccff_tail));

	sb_1__1_ sb_14__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__262_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__256_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__261_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__237_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__203_ccff_tail),
		.chany_top_out(sb_1__1__222_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__222_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__222_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__222_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__222_ccff_tail));

	sb_1__1_ sb_14__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__263_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__257_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__262_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__238_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__242_ccff_tail),
		.chany_top_out(sb_1__1__223_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__223_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__223_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__223_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__223_ccff_tail));

	sb_1__1_ sb_14__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__264_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__258_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__263_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__239_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__205_ccff_tail),
		.chany_top_out(sb_1__1__224_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__224_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__224_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__224_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__224_ccff_tail));

	sb_1__1_ sb_14__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__265_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__259_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__264_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__240_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__244_ccff_tail),
		.chany_top_out(sb_1__1__225_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__225_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__225_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__225_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__225_ccff_tail));

	sb_1__1_ sb_14__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__266_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__260_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__265_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__241_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__207_ccff_tail),
		.chany_top_out(sb_1__1__226_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__226_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__226_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__226_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__226_ccff_tail));

	sb_1__1_ sb_14__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__267_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__261_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__266_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__242_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__246_ccff_tail),
		.chany_top_out(sb_1__1__227_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__227_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__227_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__227_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__227_ccff_tail));

	sb_1__1_ sb_14__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__268_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__262_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__267_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__243_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__209_ccff_tail),
		.chany_top_out(sb_1__1__228_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__228_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__228_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__228_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__228_ccff_tail));

	sb_1__1_ sb_14__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__269_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__263_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__268_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__244_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__248_ccff_tail),
		.chany_top_out(sb_1__1__229_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__229_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__229_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__229_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__229_ccff_tail));

	sb_1__1_ sb_14__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__270_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__264_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__269_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__245_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__211_ccff_tail),
		.chany_top_out(sb_1__1__230_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__230_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__230_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__230_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__230_ccff_tail));

	sb_1__1_ sb_14__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__271_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__265_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__270_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__246_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__250_ccff_tail),
		.chany_top_out(sb_1__1__231_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__231_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__231_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__231_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__231_ccff_tail));

	sb_1__1_ sb_14__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__272_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__266_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__271_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__247_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__213_ccff_tail),
		.chany_top_out(sb_1__1__232_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__232_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__232_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__232_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__232_ccff_tail));

	sb_1__1_ sb_14__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__273_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__267_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__272_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__248_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__252_ccff_tail),
		.chany_top_out(sb_1__1__233_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__233_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__233_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__233_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__233_ccff_tail));

	sb_1__1_ sb_14__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__274_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__268_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__273_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__249_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__215_ccff_tail),
		.chany_top_out(sb_1__1__234_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__234_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__234_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__234_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__234_ccff_tail));

	sb_1__1_ sb_14__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__275_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__269_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__274_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__250_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__254_ccff_tail),
		.chany_top_out(sb_1__1__235_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__235_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__235_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__235_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__235_ccff_tail));

	sb_1__1_ sb_15__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__277_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__270_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__276_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__251_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__255_ccff_tail),
		.chany_top_out(sb_1__1__236_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__236_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__236_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__236_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__236_ccff_tail));

	sb_1__1_ sb_15__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__278_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__271_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__277_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__252_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__218_ccff_tail),
		.chany_top_out(sb_1__1__237_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__237_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__237_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__237_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__237_ccff_tail));

	sb_1__1_ sb_15__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__279_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__272_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__278_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__253_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__257_ccff_tail),
		.chany_top_out(sb_1__1__238_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__238_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__238_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__238_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__238_ccff_tail));

	sb_1__1_ sb_15__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__281_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__273_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__280_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__254_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__220_ccff_tail),
		.chany_top_out(sb_1__1__239_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__239_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__239_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__239_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__239_ccff_tail));

	sb_1__1_ sb_15__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__282_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__274_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__281_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__255_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__259_ccff_tail),
		.chany_top_out(sb_1__1__240_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__240_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__240_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__240_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__240_ccff_tail));

	sb_1__1_ sb_15__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__283_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__275_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__282_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__256_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__222_ccff_tail),
		.chany_top_out(sb_1__1__241_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__241_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__241_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__241_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__241_ccff_tail));

	sb_1__1_ sb_15__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__284_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__276_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__283_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__257_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__261_ccff_tail),
		.chany_top_out(sb_1__1__242_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__242_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__242_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__242_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__242_ccff_tail));

	sb_1__1_ sb_15__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__285_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__277_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__284_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__258_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__224_ccff_tail),
		.chany_top_out(sb_1__1__243_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__243_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__243_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__243_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__243_ccff_tail));

	sb_1__1_ sb_15__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__286_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__278_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__285_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__259_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__263_ccff_tail),
		.chany_top_out(sb_1__1__244_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__244_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__244_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__244_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__244_ccff_tail));

	sb_1__1_ sb_15__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__287_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__279_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__286_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__260_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__226_ccff_tail),
		.chany_top_out(sb_1__1__245_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__245_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__245_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__245_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__245_ccff_tail));

	sb_1__1_ sb_15__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__288_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__280_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__287_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__261_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__265_ccff_tail),
		.chany_top_out(sb_1__1__246_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__246_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__246_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__246_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__246_ccff_tail));

	sb_1__1_ sb_15__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__289_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__281_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__288_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__262_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__228_ccff_tail),
		.chany_top_out(sb_1__1__247_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__247_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__247_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__247_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__247_ccff_tail));

	sb_1__1_ sb_15__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__290_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__282_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__289_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__263_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__267_ccff_tail),
		.chany_top_out(sb_1__1__248_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__248_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__248_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__248_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__248_ccff_tail));

	sb_1__1_ sb_15__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__291_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__283_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__290_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__264_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__230_ccff_tail),
		.chany_top_out(sb_1__1__249_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__249_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__249_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__249_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__249_ccff_tail));

	sb_1__1_ sb_15__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__292_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__284_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__291_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__265_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__269_ccff_tail),
		.chany_top_out(sb_1__1__250_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__250_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__250_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__250_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__250_ccff_tail));

	sb_1__1_ sb_15__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__293_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__285_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__292_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__266_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__232_ccff_tail),
		.chany_top_out(sb_1__1__251_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__251_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__251_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__251_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__251_ccff_tail));

	sb_1__1_ sb_15__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__294_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__286_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__293_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__267_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__271_ccff_tail),
		.chany_top_out(sb_1__1__252_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__252_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__252_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__252_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__252_ccff_tail));

	sb_1__1_ sb_15__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__295_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__287_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__294_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__268_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__234_ccff_tail),
		.chany_top_out(sb_1__1__253_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__253_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__253_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__253_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__253_ccff_tail));

	sb_1__1_ sb_15__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__296_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__288_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__295_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__269_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__273_ccff_tail),
		.chany_top_out(sb_1__1__254_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__254_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__254_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__254_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__254_ccff_tail));

	sb_1__1_ sb_16__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__298_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__289_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__297_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__270_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__274_ccff_tail),
		.chany_top_out(sb_1__1__255_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__255_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__255_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__255_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__255_ccff_tail));

	sb_1__1_ sb_16__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__299_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__290_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__298_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__271_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__237_ccff_tail),
		.chany_top_out(sb_1__1__256_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__256_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__256_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__256_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__256_ccff_tail));

	sb_1__1_ sb_16__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__300_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__291_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__299_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__272_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__276_ccff_tail),
		.chany_top_out(sb_1__1__257_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__257_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__257_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__257_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__257_ccff_tail));

	sb_1__1_ sb_16__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__302_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__292_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__301_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__273_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__239_ccff_tail),
		.chany_top_out(sb_1__1__258_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__258_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__258_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__258_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__258_ccff_tail));

	sb_1__1_ sb_16__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__303_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__293_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__302_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__274_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__278_ccff_tail),
		.chany_top_out(sb_1__1__259_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__259_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__259_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__259_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__259_ccff_tail));

	sb_1__1_ sb_16__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__304_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__294_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__303_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__275_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__241_ccff_tail),
		.chany_top_out(sb_1__1__260_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__260_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__260_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__260_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__260_ccff_tail));

	sb_1__1_ sb_16__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__305_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__295_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__304_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__276_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__280_ccff_tail),
		.chany_top_out(sb_1__1__261_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__261_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__261_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__261_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__261_ccff_tail));

	sb_1__1_ sb_16__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__306_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__296_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__305_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__277_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__243_ccff_tail),
		.chany_top_out(sb_1__1__262_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__262_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__262_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__262_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__262_ccff_tail));

	sb_1__1_ sb_16__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__307_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__297_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__306_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__278_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__282_ccff_tail),
		.chany_top_out(sb_1__1__263_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__263_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__263_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__263_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__263_ccff_tail));

	sb_1__1_ sb_16__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__308_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__298_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__307_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__279_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__245_ccff_tail),
		.chany_top_out(sb_1__1__264_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__264_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__264_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__264_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__264_ccff_tail));

	sb_1__1_ sb_16__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__309_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__299_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__308_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__280_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__284_ccff_tail),
		.chany_top_out(sb_1__1__265_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__265_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__265_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__265_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__265_ccff_tail));

	sb_1__1_ sb_16__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__310_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__300_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__309_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__281_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__247_ccff_tail),
		.chany_top_out(sb_1__1__266_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__266_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__266_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__266_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__266_ccff_tail));

	sb_1__1_ sb_16__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__311_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__301_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__310_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__282_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__286_ccff_tail),
		.chany_top_out(sb_1__1__267_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__267_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__267_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__267_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__267_ccff_tail));

	sb_1__1_ sb_16__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__312_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__302_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__311_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__283_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__249_ccff_tail),
		.chany_top_out(sb_1__1__268_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__268_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__268_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__268_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__268_ccff_tail));

	sb_1__1_ sb_16__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__313_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__303_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__312_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__284_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__288_ccff_tail),
		.chany_top_out(sb_1__1__269_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__269_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__269_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__269_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__269_ccff_tail));

	sb_1__1_ sb_16__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__314_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__304_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__313_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__285_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__251_ccff_tail),
		.chany_top_out(sb_1__1__270_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__270_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__270_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__270_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__270_ccff_tail));

	sb_1__1_ sb_16__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__315_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__305_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__314_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__286_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__290_ccff_tail),
		.chany_top_out(sb_1__1__271_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__271_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__271_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__271_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__271_ccff_tail));

	sb_1__1_ sb_16__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__316_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__306_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__315_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__287_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__253_ccff_tail),
		.chany_top_out(sb_1__1__272_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__272_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__272_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__272_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__272_ccff_tail));

	sb_1__1_ sb_16__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__317_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__307_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__316_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__288_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__292_ccff_tail),
		.chany_top_out(sb_1__1__273_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__273_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__273_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__273_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__273_ccff_tail));

	sb_1__1_ sb_17__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__319_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__308_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__318_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__289_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__293_ccff_tail),
		.chany_top_out(sb_1__1__274_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__274_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__274_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__274_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__274_ccff_tail));

	sb_1__1_ sb_17__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__320_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__309_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__319_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__290_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__256_ccff_tail),
		.chany_top_out(sb_1__1__275_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__275_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__275_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__275_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__275_ccff_tail));

	sb_1__1_ sb_17__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__321_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__310_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__320_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__291_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__295_ccff_tail),
		.chany_top_out(sb_1__1__276_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__276_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__276_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__276_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__276_ccff_tail));

	sb_1__1_ sb_17__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__323_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__311_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__322_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__292_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__258_ccff_tail),
		.chany_top_out(sb_1__1__277_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__277_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__277_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__277_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__277_ccff_tail));

	sb_1__1_ sb_17__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__324_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__312_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__323_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__293_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__297_ccff_tail),
		.chany_top_out(sb_1__1__278_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__278_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__278_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__278_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__278_ccff_tail));

	sb_1__1_ sb_17__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__325_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__313_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__324_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__294_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__260_ccff_tail),
		.chany_top_out(sb_1__1__279_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__279_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__279_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__279_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__279_ccff_tail));

	sb_1__1_ sb_17__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__326_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__314_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__325_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__295_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__299_ccff_tail),
		.chany_top_out(sb_1__1__280_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__280_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__280_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__280_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__280_ccff_tail));

	sb_1__1_ sb_17__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__327_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__315_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__326_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__296_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__262_ccff_tail),
		.chany_top_out(sb_1__1__281_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__281_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__281_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__281_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__281_ccff_tail));

	sb_1__1_ sb_17__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__328_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__316_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__327_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__297_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__301_ccff_tail),
		.chany_top_out(sb_1__1__282_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__282_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__282_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__282_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__282_ccff_tail));

	sb_1__1_ sb_17__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__329_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__317_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__328_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__298_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__264_ccff_tail),
		.chany_top_out(sb_1__1__283_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__283_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__283_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__283_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__283_ccff_tail));

	sb_1__1_ sb_17__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__330_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__318_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__329_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__299_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__303_ccff_tail),
		.chany_top_out(sb_1__1__284_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__284_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__284_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__284_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__284_ccff_tail));

	sb_1__1_ sb_17__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__331_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__319_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__330_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__300_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__266_ccff_tail),
		.chany_top_out(sb_1__1__285_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__285_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__285_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__285_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__285_ccff_tail));

	sb_1__1_ sb_17__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__332_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__320_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__331_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__301_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__305_ccff_tail),
		.chany_top_out(sb_1__1__286_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__286_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__286_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__286_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__286_ccff_tail));

	sb_1__1_ sb_17__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__333_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__321_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__332_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__302_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__268_ccff_tail),
		.chany_top_out(sb_1__1__287_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__287_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__287_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__287_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__287_ccff_tail));

	sb_1__1_ sb_17__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__334_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__322_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__333_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__303_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__307_ccff_tail),
		.chany_top_out(sb_1__1__288_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__288_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__288_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__288_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__288_ccff_tail));

	sb_1__1_ sb_17__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__335_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__323_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__334_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__304_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__270_ccff_tail),
		.chany_top_out(sb_1__1__289_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__289_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__289_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__289_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__289_ccff_tail));

	sb_1__1_ sb_17__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__336_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__324_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__335_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__305_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__309_ccff_tail),
		.chany_top_out(sb_1__1__290_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__290_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__290_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__290_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__290_ccff_tail));

	sb_1__1_ sb_17__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__337_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__325_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__336_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__306_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__272_ccff_tail),
		.chany_top_out(sb_1__1__291_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__291_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__291_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__291_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__291_ccff_tail));

	sb_1__1_ sb_17__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__338_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__326_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__337_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__307_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__311_ccff_tail),
		.chany_top_out(sb_1__1__292_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__292_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__292_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__292_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__292_ccff_tail));

	sb_1__1_ sb_18__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__340_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__327_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__339_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__308_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__312_ccff_tail),
		.chany_top_out(sb_1__1__293_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__293_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__293_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__293_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__293_ccff_tail));

	sb_1__1_ sb_18__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__341_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__328_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__340_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__309_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__275_ccff_tail),
		.chany_top_out(sb_1__1__294_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__294_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__294_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__294_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__294_ccff_tail));

	sb_1__1_ sb_18__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__342_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__329_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__341_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__310_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__314_ccff_tail),
		.chany_top_out(sb_1__1__295_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__295_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__295_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__295_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__295_ccff_tail));

	sb_1__1_ sb_18__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__344_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__330_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__343_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__311_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__277_ccff_tail),
		.chany_top_out(sb_1__1__296_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__296_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__296_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__296_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__296_ccff_tail));

	sb_1__1_ sb_18__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__345_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__331_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__344_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__312_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__316_ccff_tail),
		.chany_top_out(sb_1__1__297_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__297_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__297_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__297_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__297_ccff_tail));

	sb_1__1_ sb_18__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__346_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__332_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__345_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__313_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__279_ccff_tail),
		.chany_top_out(sb_1__1__298_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__298_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__298_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__298_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__298_ccff_tail));

	sb_1__1_ sb_18__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__347_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__333_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__346_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__314_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__318_ccff_tail),
		.chany_top_out(sb_1__1__299_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__299_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__299_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__299_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__299_ccff_tail));

	sb_1__1_ sb_18__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__348_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__334_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__347_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__315_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__281_ccff_tail),
		.chany_top_out(sb_1__1__300_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__300_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__300_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__300_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__300_ccff_tail));

	sb_1__1_ sb_18__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__349_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__335_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__348_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__316_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__320_ccff_tail),
		.chany_top_out(sb_1__1__301_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__301_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__301_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__301_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__301_ccff_tail));

	sb_1__1_ sb_18__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__350_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__336_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__349_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__317_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__283_ccff_tail),
		.chany_top_out(sb_1__1__302_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__302_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__302_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__302_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__302_ccff_tail));

	sb_1__1_ sb_18__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__351_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__337_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__350_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__318_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__322_ccff_tail),
		.chany_top_out(sb_1__1__303_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__303_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__303_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__303_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__303_ccff_tail));

	sb_1__1_ sb_18__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__352_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__338_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__351_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__319_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__285_ccff_tail),
		.chany_top_out(sb_1__1__304_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__304_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__304_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__304_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__304_ccff_tail));

	sb_1__1_ sb_18__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__353_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__339_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__352_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__320_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__324_ccff_tail),
		.chany_top_out(sb_1__1__305_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__305_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__305_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__305_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__305_ccff_tail));

	sb_1__1_ sb_18__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__354_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__340_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__353_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__321_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__287_ccff_tail),
		.chany_top_out(sb_1__1__306_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__306_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__306_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__306_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__306_ccff_tail));

	sb_1__1_ sb_18__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__355_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__341_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__354_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__322_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__326_ccff_tail),
		.chany_top_out(sb_1__1__307_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__307_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__307_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__307_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__307_ccff_tail));

	sb_1__1_ sb_18__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__356_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__342_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__355_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__323_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__289_ccff_tail),
		.chany_top_out(sb_1__1__308_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__308_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__308_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__308_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__308_ccff_tail));

	sb_1__1_ sb_18__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__357_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__343_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__356_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__324_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__328_ccff_tail),
		.chany_top_out(sb_1__1__309_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__309_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__309_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__309_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__309_ccff_tail));

	sb_1__1_ sb_18__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__358_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__344_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__357_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__325_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__291_ccff_tail),
		.chany_top_out(sb_1__1__310_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__310_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__310_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__310_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__310_ccff_tail));

	sb_1__1_ sb_18__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__359_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__345_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__358_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__326_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__330_ccff_tail),
		.chany_top_out(sb_1__1__311_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__311_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__311_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__311_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__311_ccff_tail));

	sb_1__1_ sb_19__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__361_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__346_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__360_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__327_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__331_ccff_tail),
		.chany_top_out(sb_1__1__312_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__312_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__312_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__312_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__312_ccff_tail));

	sb_1__1_ sb_19__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__362_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__347_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__361_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__328_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__294_ccff_tail),
		.chany_top_out(sb_1__1__313_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__313_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__313_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__313_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__313_ccff_tail));

	sb_1__1_ sb_19__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__363_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__348_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__362_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__329_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__333_ccff_tail),
		.chany_top_out(sb_1__1__314_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__314_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__314_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__314_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__314_ccff_tail));

	sb_1__1_ sb_19__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__365_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__349_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__364_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__330_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__296_ccff_tail),
		.chany_top_out(sb_1__1__315_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__315_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__315_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__315_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__315_ccff_tail));

	sb_1__1_ sb_19__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__366_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__350_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__365_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__331_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__335_ccff_tail),
		.chany_top_out(sb_1__1__316_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__316_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__316_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__316_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__316_ccff_tail));

	sb_1__1_ sb_19__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__367_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__351_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__366_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__332_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__298_ccff_tail),
		.chany_top_out(sb_1__1__317_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__317_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__317_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__317_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__317_ccff_tail));

	sb_1__1_ sb_19__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__368_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__352_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__367_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__333_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__337_ccff_tail),
		.chany_top_out(sb_1__1__318_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__318_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__318_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__318_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__318_ccff_tail));

	sb_1__1_ sb_19__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__369_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__353_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__368_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__334_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__300_ccff_tail),
		.chany_top_out(sb_1__1__319_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__319_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__319_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__319_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__319_ccff_tail));

	sb_1__1_ sb_19__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__370_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__354_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__369_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__335_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__339_ccff_tail),
		.chany_top_out(sb_1__1__320_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__320_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__320_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__320_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__320_ccff_tail));

	sb_1__1_ sb_19__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__371_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__355_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__370_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__336_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__302_ccff_tail),
		.chany_top_out(sb_1__1__321_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__321_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__321_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__321_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__321_ccff_tail));

	sb_1__1_ sb_19__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__372_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__356_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__371_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__337_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__341_ccff_tail),
		.chany_top_out(sb_1__1__322_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__322_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__322_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__322_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__322_ccff_tail));

	sb_1__1_ sb_19__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__373_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__357_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__372_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__338_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__304_ccff_tail),
		.chany_top_out(sb_1__1__323_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__323_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__323_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__323_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__323_ccff_tail));

	sb_1__1_ sb_19__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__374_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__358_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__373_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__339_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__343_ccff_tail),
		.chany_top_out(sb_1__1__324_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__324_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__324_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__324_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__324_ccff_tail));

	sb_1__1_ sb_19__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__375_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__359_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__374_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__340_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__306_ccff_tail),
		.chany_top_out(sb_1__1__325_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__325_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__325_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__325_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__325_ccff_tail));

	sb_1__1_ sb_19__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__376_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__360_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__375_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__341_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__345_ccff_tail),
		.chany_top_out(sb_1__1__326_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__326_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__326_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__326_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__326_ccff_tail));

	sb_1__1_ sb_19__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__377_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__361_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__376_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__342_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__308_ccff_tail),
		.chany_top_out(sb_1__1__327_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__327_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__327_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__327_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__327_ccff_tail));

	sb_1__1_ sb_19__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__378_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__362_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__377_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__343_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__347_ccff_tail),
		.chany_top_out(sb_1__1__328_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__328_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__328_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__328_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__328_ccff_tail));

	sb_1__1_ sb_19__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__379_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__363_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__378_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__344_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__310_ccff_tail),
		.chany_top_out(sb_1__1__329_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__329_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__329_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__329_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__329_ccff_tail));

	sb_1__1_ sb_19__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__380_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__364_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__379_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__345_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__349_ccff_tail),
		.chany_top_out(sb_1__1__330_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__330_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__330_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__330_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__330_ccff_tail));

	sb_1__1_ sb_20__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__382_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__365_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__381_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__346_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__350_ccff_tail),
		.chany_top_out(sb_1__1__331_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__331_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__331_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__331_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__331_ccff_tail));

	sb_1__1_ sb_20__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__383_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__366_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__382_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__347_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__313_ccff_tail),
		.chany_top_out(sb_1__1__332_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__332_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__332_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__332_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__332_ccff_tail));

	sb_1__1_ sb_20__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__384_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__367_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__383_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__348_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__352_ccff_tail),
		.chany_top_out(sb_1__1__333_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__333_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__333_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__333_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__333_ccff_tail));

	sb_1__1_ sb_20__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__386_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__368_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__385_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__349_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__315_ccff_tail),
		.chany_top_out(sb_1__1__334_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__334_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__334_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__334_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__334_ccff_tail));

	sb_1__1_ sb_20__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__387_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__369_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__386_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__350_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__354_ccff_tail),
		.chany_top_out(sb_1__1__335_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__335_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__335_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__335_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__335_ccff_tail));

	sb_1__1_ sb_20__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__388_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__370_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__387_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__351_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__317_ccff_tail),
		.chany_top_out(sb_1__1__336_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__336_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__336_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__336_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__336_ccff_tail));

	sb_1__1_ sb_20__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__389_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__371_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__388_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__352_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__356_ccff_tail),
		.chany_top_out(sb_1__1__337_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__337_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__337_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__337_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__337_ccff_tail));

	sb_1__1_ sb_20__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__390_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__372_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__389_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__353_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__319_ccff_tail),
		.chany_top_out(sb_1__1__338_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__338_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__338_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__338_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__338_ccff_tail));

	sb_1__1_ sb_20__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__391_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__373_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__390_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__354_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__358_ccff_tail),
		.chany_top_out(sb_1__1__339_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__339_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__339_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__339_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__339_ccff_tail));

	sb_1__1_ sb_20__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__392_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__374_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__391_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__355_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__321_ccff_tail),
		.chany_top_out(sb_1__1__340_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__340_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__340_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__340_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__340_ccff_tail));

	sb_1__1_ sb_20__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__393_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__375_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__392_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__356_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__360_ccff_tail),
		.chany_top_out(sb_1__1__341_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__341_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__341_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__341_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__341_ccff_tail));

	sb_1__1_ sb_20__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__394_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__376_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__393_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__357_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__323_ccff_tail),
		.chany_top_out(sb_1__1__342_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__342_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__342_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__342_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__342_ccff_tail));

	sb_1__1_ sb_20__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__395_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__377_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__394_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__358_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__362_ccff_tail),
		.chany_top_out(sb_1__1__343_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__343_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__343_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__343_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__343_ccff_tail));

	sb_1__1_ sb_20__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__396_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__378_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__395_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__359_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__325_ccff_tail),
		.chany_top_out(sb_1__1__344_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__344_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__344_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__344_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__344_ccff_tail));

	sb_1__1_ sb_20__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__397_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__379_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__396_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__360_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__364_ccff_tail),
		.chany_top_out(sb_1__1__345_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__345_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__345_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__345_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__345_ccff_tail));

	sb_1__1_ sb_20__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__398_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__380_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__397_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__361_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__327_ccff_tail),
		.chany_top_out(sb_1__1__346_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__346_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__346_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__346_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__346_ccff_tail));

	sb_1__1_ sb_20__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__399_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__381_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__398_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__362_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__366_ccff_tail),
		.chany_top_out(sb_1__1__347_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__347_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__347_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__347_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__347_ccff_tail));

	sb_1__1_ sb_20__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__400_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__382_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__399_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__363_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__329_ccff_tail),
		.chany_top_out(sb_1__1__348_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__348_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__348_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__348_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__348_ccff_tail));

	sb_1__1_ sb_20__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__401_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__383_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__400_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__364_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__368_ccff_tail),
		.chany_top_out(sb_1__1__349_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__349_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__349_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__349_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__349_ccff_tail));

	sb_1__1_ sb_21__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__403_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__384_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__402_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__365_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__1_ccff_tail),
		.chany_top_out(sb_1__1__350_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__350_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__350_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__350_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__350_ccff_tail));

	sb_1__1_ sb_21__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__404_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__385_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__403_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__366_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__332_ccff_tail),
		.chany_top_out(sb_1__1__351_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__351_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__351_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__351_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__351_ccff_tail));

	sb_1__1_ sb_21__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__405_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__386_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__404_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__367_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__3_ccff_tail),
		.chany_top_out(sb_1__1__352_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__352_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__352_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__352_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__352_ccff_tail));

	sb_1__1_ sb_21__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__407_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__387_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__406_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__368_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__334_ccff_tail),
		.chany_top_out(sb_1__1__353_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__353_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__353_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__353_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__353_ccff_tail));

	sb_1__1_ sb_21__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__408_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__388_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__407_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__369_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__6_ccff_tail),
		.chany_top_out(sb_1__1__354_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__354_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__354_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__354_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__354_ccff_tail));

	sb_1__1_ sb_21__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__409_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__389_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__408_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__370_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__336_ccff_tail),
		.chany_top_out(sb_1__1__355_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__355_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__355_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__355_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__355_ccff_tail));

	sb_1__1_ sb_21__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__410_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__390_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__409_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__371_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__8_ccff_tail),
		.chany_top_out(sb_1__1__356_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__356_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__356_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__356_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__356_ccff_tail));

	sb_1__1_ sb_21__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__411_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__391_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__410_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__372_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__338_ccff_tail),
		.chany_top_out(sb_1__1__357_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__357_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__357_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__357_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__357_ccff_tail));

	sb_1__1_ sb_21__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__412_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__392_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__411_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__373_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__10_ccff_tail),
		.chany_top_out(sb_1__1__358_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__358_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__358_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__358_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__358_ccff_tail));

	sb_1__1_ sb_21__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__413_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__393_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__412_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__374_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__340_ccff_tail),
		.chany_top_out(sb_1__1__359_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__359_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__359_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__359_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__359_ccff_tail));

	sb_1__1_ sb_21__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__414_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__394_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__413_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__375_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__12_ccff_tail),
		.chany_top_out(sb_1__1__360_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__360_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__360_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__360_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__360_ccff_tail));

	sb_1__1_ sb_21__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__415_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__395_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__414_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__376_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__342_ccff_tail),
		.chany_top_out(sb_1__1__361_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__361_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__361_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__361_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__361_ccff_tail));

	sb_1__1_ sb_21__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__416_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__396_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__415_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__377_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__14_ccff_tail),
		.chany_top_out(sb_1__1__362_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__362_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__362_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__362_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__362_ccff_tail));

	sb_1__1_ sb_21__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__417_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__397_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__416_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__378_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__344_ccff_tail),
		.chany_top_out(sb_1__1__363_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__363_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__363_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__363_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__363_ccff_tail));

	sb_1__1_ sb_21__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__418_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__398_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__417_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__379_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__16_ccff_tail),
		.chany_top_out(sb_1__1__364_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__364_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__364_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__364_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__364_ccff_tail));

	sb_1__1_ sb_21__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__419_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__399_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__418_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__380_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__346_ccff_tail),
		.chany_top_out(sb_1__1__365_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__365_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__365_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__365_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__365_ccff_tail));

	sb_1__1_ sb_21__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__420_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__400_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__419_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__381_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__18_ccff_tail),
		.chany_top_out(sb_1__1__366_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__366_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__366_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__366_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__366_ccff_tail));

	sb_1__1_ sb_21__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__421_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__401_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__420_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__382_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__348_ccff_tail),
		.chany_top_out(sb_1__1__367_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__367_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__367_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__367_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__367_ccff_tail));

	sb_1__1_ sb_21__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__422_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__402_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__421_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__383_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__20_ccff_tail),
		.chany_top_out(sb_1__1__368_chany_top_out[0:228]),
		.chanx_right_out(sb_1__1__368_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__1__368_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__1__368_chanx_left_out[0:228]),
		.ccff_tail(sb_1__1__368_ccff_tail));

	sb_1__4_ sb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__0_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__1_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__0_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chany_top_out(sb_1__4__0_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__0_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__0_ccff_tail));

	sb_1__4_ sb_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__1_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__2_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__1_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__4__1_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__1_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__1_ccff_tail));

	sb_1__4_ sb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__2_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__3_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__2_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__4__2_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__2_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__2_ccff_tail));

	sb_1__4_ sb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__3_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__4_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__60_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__3_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__4__3_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__3_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__3_ccff_tail));

	sb_1__4_ sb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__4_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__5_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__80_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__4_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__4__4_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__4_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__4_ccff_tail));

	sb_1__4_ sb_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__5_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__6_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__98_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__5_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__4__5_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__5_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__5_ccff_tail));

	sb_1__4_ sb_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__6_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__7_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__117_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__6_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__4__6_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__6_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__6_ccff_tail));

	sb_1__4_ sb_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__7_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__8_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__137_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__7_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__4__7_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__7_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__7_ccff_tail));

	sb_1__4_ sb_9__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__8_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__9_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__155_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__8_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__4__8_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__8_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__8_ccff_tail));

	sb_1__4_ sb_10__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__9_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__10_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__174_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__9_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__4__9_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__9_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__9_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__9_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__9_ccff_tail));

	sb_1__4_ sb_11__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__10_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__11_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__195_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__10_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__4__10_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__10_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__10_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__10_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__10_ccff_tail));

	sb_1__4_ sb_12__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__11_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__12_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__216_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__11_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__4__11_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__11_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__11_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__11_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__11_ccff_tail));

	sb_1__4_ sb_13__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__12_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__13_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__237_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__12_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__4__12_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__12_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__12_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__12_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__12_ccff_tail));

	sb_1__4_ sb_14__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__13_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__14_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__258_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__13_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__4__13_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__13_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__13_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__13_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__13_ccff_tail));

	sb_1__4_ sb_15__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__14_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__15_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__279_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__14_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__4__14_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__14_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__14_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__14_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__14_ccff_tail));

	sb_1__4_ sb_16__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__15_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__16_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__300_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__15_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__4__15_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__15_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__15_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__15_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__15_ccff_tail));

	sb_1__4_ sb_17__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__16_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__17_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__321_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__16_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__4__16_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__16_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__16_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__16_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__16_ccff_tail));

	sb_1__4_ sb_18__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__17_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__18_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__342_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__17_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__4__17_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__17_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__17_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__17_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__17_ccff_tail));

	sb_1__4_ sb_19__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__18_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__19_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__363_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__18_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_1__4__18_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__18_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__18_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__18_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__18_ccff_tail));

	sb_1__4_ sb_20__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__19_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__20_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__384_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__19_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__4__19_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__19_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__19_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__19_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__19_ccff_tail));

	sb_1__4_ sb_21__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__5__20_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__4__21_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.chany_bottom_in(cby_1__1__405_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__4__20_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_1__4__20_chany_top_out[0:228]),
		.chanx_right_out(sb_1__4__20_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__4__20_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__4__20_chanx_left_out[0:228]),
		.ccff_tail(sb_1__4__20_ccff_tail));

	sb_1__5_ sb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__1_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__0_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__0_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_2__3__1_ccff_tail),
		.chany_top_out(sb_1__5__0_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__0_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__0_ccff_tail));

	sb_1__5_ sb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__61_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__3_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__3_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__2_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_2__3__4_ccff_tail),
		.chany_top_out(sb_1__5__1_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__1_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__1_ccff_tail));

	sb_1__5_ sb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__118_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__5_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__6_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__4_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_2__3__7_ccff_tail),
		.chany_top_out(sb_1__5__2_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__2_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__2_ccff_tail));

	sb_1__5_ sb_10__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__175_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__7_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__9_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__6_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__7_ccff_tail),
		.chany_top_out(sb_1__5__3_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__3_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__3_ccff_tail));

	sb_1__5_ sb_11__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__196_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__8_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__10_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__7_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__8_ccff_tail),
		.chany_top_out(sb_1__5__4_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__4_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__4_ccff_tail));

	sb_1__5_ sb_12__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__217_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__9_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__11_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__8_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__9_ccff_tail),
		.chany_top_out(sb_1__5__5_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__5_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__5_ccff_tail));

	sb_1__5_ sb_13__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__238_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__10_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__12_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__9_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__10_ccff_tail),
		.chany_top_out(sb_1__5__6_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__6_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__6_ccff_tail));

	sb_1__5_ sb_14__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__259_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__11_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__13_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__10_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__11_ccff_tail),
		.chany_top_out(sb_1__5__7_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__7_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__7_ccff_tail));

	sb_1__5_ sb_15__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__280_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__12_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__14_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__11_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__12_ccff_tail),
		.chany_top_out(sb_1__5__8_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__8_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__8_ccff_tail));

	sb_1__5_ sb_16__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__301_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__13_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__15_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__12_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__13_ccff_tail),
		.chany_top_out(sb_1__5__9_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__9_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__9_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__9_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__9_ccff_tail));

	sb_1__5_ sb_17__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__322_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__14_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__16_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__13_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__14_ccff_tail),
		.chany_top_out(sb_1__5__10_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__10_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__10_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__10_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__10_ccff_tail));

	sb_1__5_ sb_18__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__343_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__15_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__17_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__14_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__15_ccff_tail),
		.chany_top_out(sb_1__5__11_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__11_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__11_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__11_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__11_ccff_tail));

	sb_1__5_ sb_19__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__364_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__16_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__18_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__15_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__16_ccff_tail),
		.chany_top_out(sb_1__5__12_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__12_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__12_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__12_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__12_ccff_tail));

	sb_1__5_ sb_20__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__385_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__17_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__19_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__16_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__17_ccff_tail),
		.chany_top_out(sb_1__5__13_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__13_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__13_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__13_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__13_ccff_tail));

	sb_1__5_ sb_21__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__406_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__5__18_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__20_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__17_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_22__1__4_ccff_tail),
		.chany_top_out(sb_1__5__14_chany_top_out[0:228]),
		.chanx_right_out(sb_1__5__14_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__5__14_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__5__14_chanx_left_out[0:228]),
		.ccff_tail(sb_1__5__14_ccff_tail));

	sb_1__22_ sb_1__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__1_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__0_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__22__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__0_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__0_ccff_tail));

	sb_1__22_ sb_2__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__2_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__1_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__22__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__1_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__1_ccff_tail));

	sb_1__22_ sb_3__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__3_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__56_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__2_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chanx_right_out(sb_1__22__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__2_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__2_ccff_tail));

	sb_1__22_ sb_4__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__4_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__77_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__3_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_4_ccff_tail),
		.chanx_right_out(sb_1__22__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__3_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__3_ccff_tail));

	sb_1__22_ sb_5__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__5_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__95_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__4_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_5_ccff_tail),
		.chanx_right_out(sb_1__22__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__4_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__4_ccff_tail));

	sb_1__22_ sb_6__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__6_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__113_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__5_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_6_ccff_tail),
		.chanx_right_out(sb_1__22__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__5_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__5_ccff_tail));

	sb_1__22_ sb_7__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__7_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__134_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__6_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_7_ccff_tail),
		.chanx_right_out(sb_1__22__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__6_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__6_ccff_tail));

	sb_1__22_ sb_8__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__8_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__152_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__7_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_8_ccff_tail),
		.chanx_right_out(sb_1__22__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__7_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__7_ccff_tail));

	sb_1__22_ sb_9__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__9_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__170_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__8_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_9_ccff_tail),
		.chanx_right_out(sb_1__22__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__8_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__8_ccff_tail));

	sb_1__22_ sb_10__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__10_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__191_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__9_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_10_ccff_tail),
		.chanx_right_out(sb_1__22__9_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__9_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__9_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__9_ccff_tail));

	sb_1__22_ sb_11__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__11_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__212_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__10_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_11_ccff_tail),
		.chanx_right_out(sb_1__22__10_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__10_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__10_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__10_ccff_tail));

	sb_1__22_ sb_12__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__12_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__233_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__11_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_12_ccff_tail),
		.chanx_right_out(sb_1__22__11_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__11_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__11_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__11_ccff_tail));

	sb_1__22_ sb_13__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__13_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__254_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__12_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_13_ccff_tail),
		.chanx_right_out(sb_1__22__12_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__12_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__12_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__12_ccff_tail));

	sb_1__22_ sb_14__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__14_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__275_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__13_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_14_ccff_tail),
		.chanx_right_out(sb_1__22__13_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__13_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__13_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__13_ccff_tail));

	sb_1__22_ sb_15__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__15_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__296_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__14_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_15_ccff_tail),
		.chanx_right_out(sb_1__22__14_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__14_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__14_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__14_ccff_tail));

	sb_1__22_ sb_16__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__16_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__317_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__15_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_16_ccff_tail),
		.chanx_right_out(sb_1__22__15_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__15_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__15_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__15_ccff_tail));

	sb_1__22_ sb_17__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__17_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__338_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__16_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_17_ccff_tail),
		.chanx_right_out(sb_1__22__16_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__16_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__16_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__16_ccff_tail));

	sb_1__22_ sb_18__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__18_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__359_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__17_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_18_ccff_tail),
		.chanx_right_out(sb_1__22__17_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__17_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__17_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__17_ccff_tail));

	sb_1__22_ sb_19__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__19_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__380_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__18_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_19_ccff_tail),
		.chanx_right_out(sb_1__22__18_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__18_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__18_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__18_ccff_tail));

	sb_1__22_ sb_20__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__20_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__401_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__19_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_20_ccff_tail),
		.chanx_right_out(sb_1__22__19_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__19_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__19_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__19_ccff_tail));

	sb_1__22_ sb_21__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__22__21_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__1__422_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__22__20_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_20_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_21_ccff_tail),
		.chanx_right_out(sb_1__22__20_chanx_right_out[0:228]),
		.chany_bottom_out(sb_1__22__20_chany_bottom_out[0:228]),
		.chanx_left_out(sb_1__22__20_chanx_left_out[0:228]),
		.ccff_tail(sb_1__22__20_ccff_tail));

	sb_2__2_ sb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__0_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__0_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__20_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chany_top_out(sb_2__2__0_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__0_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__0_ccff_tail));

	sb_2__2_ sb_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__2_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__1_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__24_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chany_top_out(sb_2__2__1_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__1_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__1_ccff_tail));

	sb_2__2_ sb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__3_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__2_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__79_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__72_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__48_ccff_tail),
		.chany_top_out(sb_2__2__2_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__2_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__2_ccff_tail));

	sb_2__2_ sb_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__5_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__3_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__82_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__76_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__52_ccff_tail),
		.chany_top_out(sb_2__2__3_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__3_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__3_ccff_tail));

	sb_2__2_ sb_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__6_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__4_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__136_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__124_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__95_ccff_tail),
		.chany_top_out(sb_2__2__4_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__4_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__4_ccff_tail));

	sb_2__2_ sb_8__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__8_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__2__5_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.chany_bottom_in(cby_1__1__139_chany_top_out[0:228]),
		.chanx_left_in(cbx_1__1__128_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__99_ccff_tail),
		.chany_top_out(sb_2__2__5_chany_top_out[0:228]),
		.chanx_right_out(sb_2__2__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__2__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__2__5_chanx_left_out[0:228]),
		.ccff_tail(sb_2__2__5_ccff_tail));

	sb_2__3_ sb_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__23_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__0_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__0_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__21_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__0_ccff_tail),
		.chany_top_out(sb_2__3__0_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__0_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__0_ccff_tail));

	sb_2__3_ sb_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__24_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__1_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__1_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__22_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chany_top_out(sb_2__3__1_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__1_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__1_ccff_tail));

	sb_2__3_ sb_2__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__26_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__2_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__2_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_2_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__25_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__2_ccff_tail),
		.chany_top_out(sb_2__3__2_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__2_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__2_ccff_tail));

	sb_2__3_ sb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__80_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__3_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__3_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_3_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__73_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__3_ccff_tail),
		.chany_top_out(sb_2__3__3_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__3_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__3_ccff_tail));

	sb_2__3_ sb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__81_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__4_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__4_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__74_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__50_ccff_tail),
		.chany_top_out(sb_2__3__4_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__4_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__4_ccff_tail));

	sb_2__3_ sb_5__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__83_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__5_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__5_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_5_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_5_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__77_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__5_ccff_tail),
		.chany_top_out(sb_2__3__5_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__5_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__5_ccff_tail));

	sb_2__3_ sb_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__137_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__6_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__6_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_6_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_6_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__125_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__6_ccff_tail),
		.chany_top_out(sb_2__3__6_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__6_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__6_ccff_tail));

	sb_2__3_ sb_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__138_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__7_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__7_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__126_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__97_ccff_tail),
		.chany_top_out(sb_2__3__7_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__7_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__7_ccff_tail));

	sb_2__3_ sb_8__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__140_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_3__3__8_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.chany_bottom_in(cby_2__3__8_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_8_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_8_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_left_in(cbx_1__1__129_chanx_right_out[0:228]),
		.ccff_head(cbx_3__3__8_ccff_tail),
		.chany_top_out(sb_2__3__8_chany_top_out[0:228]),
		.chanx_right_out(sb_2__3__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__3__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__3__8_chanx_left_out[0:228]),
		.ccff_tail(sb_2__3__8_ccff_tail));

	sb_2__5_ sb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__1_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__5__0_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__1_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__1_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_3__3__1_ccff_tail),
		.chany_top_out(sb_2__5__0_chany_top_out[0:228]),
		.chanx_right_out(sb_2__5__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__5__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__5__0_chanx_left_out[0:228]),
		.ccff_tail(sb_2__5__0_ccff_tail));

	sb_2__5_ sb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__4_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_4_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_4_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__5__1_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__4_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__3_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_3__3__4_ccff_tail),
		.chany_top_out(sb_2__5__1_chany_top_out[0:228]),
		.chanx_right_out(sb_2__5__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__5__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__5__1_chanx_left_out[0:228]),
		.ccff_tail(sb_2__5__1_ccff_tail));

	sb_2__5_ sb_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__3__7_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_7_left_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_3_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_7_left_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chanx_right_in(cbx_3__5__2_chanx_left_out[0:228]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__7_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__5_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cby_3__3__7_ccff_tail),
		.chany_top_out(sb_2__5__2_chany_top_out[0:228]),
		.chanx_right_out(sb_2__5__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_2__5__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_2__5__2_chanx_left_out[0:228]),
		.ccff_tail(sb_2__5__2_ccff_tail));

	sb_3__2_ sb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__0_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__53_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__0_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__0_ccff_tail),
		.chany_top_out(sb_3__2__0_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__0_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__0_ccff_tail));

	sb_3__2_ sb_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__2_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__57_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__1_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__2_ccff_tail),
		.chany_top_out(sb_3__2__1_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__1_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__1_ccff_tail));

	sb_3__2_ sb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__3_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__105_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__97_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__2_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__3_ccff_tail),
		.chany_top_out(sb_3__2__2_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__2_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__2_ccff_tail));

	sb_3__2_ sb_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__5_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__109_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__100_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__3_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_5_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__5_ccff_tail),
		.chany_top_out(sb_3__2__3_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__3_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__3_ccff_tail));

	sb_3__2_ sb_9__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__6_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__157_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__154_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__4_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_6_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__6_ccff_tail),
		.chany_top_out(sb_3__2__4_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__4_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__4_ccff_tail));

	sb_3__2_ sb_9__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__8_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__1__161_chanx_left_out[0:228]),
		.chany_bottom_in(cby_1__1__157_chany_top_out[0:228]),
		.chanx_left_in(cbx_3__2__5_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_8_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.ccff_head(cby_2__3__8_ccff_tail),
		.chany_top_out(sb_3__2__5_chany_top_out[0:228]),
		.chanx_right_out(sb_3__2__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__2__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__2__5_chanx_left_out[0:228]),
		.ccff_tail(sb_3__2__5_ccff_tail));

	sb_3__3_ sb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__41_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__54_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__0_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__0_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__49_ccff_tail),
		.chany_top_out(sb_3__3__0_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__0_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__0_ccff_tail));

	sb_3__3_ sb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__42_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__55_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__1_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__1_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_2__3__1_ccff_tail),
		.chany_top_out(sb_3__3__1_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__1_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__1_ccff_tail));

	sb_3__3_ sb_3__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__44_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__58_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__2_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_2_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_2_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__2_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_2_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__53_ccff_tail),
		.chany_top_out(sb_3__3__2_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__2_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__2_ccff_tail));

	sb_3__3_ sb_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__98_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__106_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__3_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_3_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_3_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__3_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_3_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__96_ccff_tail),
		.chany_top_out(sb_3__3__3_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__3_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__3_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__3_ccff_tail));

	sb_3__3_ sb_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__99_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__107_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__4_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__4_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_4_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_4_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_2__3__4_ccff_tail),
		.chany_top_out(sb_3__3__4_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__4_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__4_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__4_ccff_tail));

	sb_3__3_ sb_6__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__101_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__110_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__5_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_5_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_5_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__5_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_5_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_5_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__100_ccff_tail),
		.chany_top_out(sb_3__3__5_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__5_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__5_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__5_ccff_tail));

	sb_3__3_ sb_9__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__155_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__158_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__6_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_6_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_6_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__6_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_6_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_6_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__143_ccff_tail),
		.chany_top_out(sb_3__3__6_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__6_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__6_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__6_ccff_tail));

	sb_3__3_ sb_9__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__156_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__159_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__7_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__7_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_7_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_7_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_2__3__7_ccff_tail),
		.chany_top_out(sb_3__3__7_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__7_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__7_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__7_ccff_tail));

	sb_3__3_ sb_9__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__158_chany_bottom_out[0:228]),
		.chanx_right_in(cbx_1__1__162_chanx_left_out[0:228]),
		.chany_bottom_in(cby_3__3__8_chany_top_out[0:228]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_8_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_8_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_left_in(cbx_3__3__8_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_8_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_8_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.ccff_head(sb_1__1__147_ccff_tail),
		.chany_top_out(sb_3__3__8_chany_top_out[0:228]),
		.chanx_right_out(sb_3__3__8_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__3__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__3__8_chanx_left_out[0:228]),
		.ccff_tail(sb_3__3__8_ccff_tail));

	sb_3__5_ sb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__1_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__5__2_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__2_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_3__5__0_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__2_ccff_tail),
		.chany_top_out(sb_3__5__0_chany_top_out[0:228]),
		.chanx_right_out(sb_3__5__0_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__5__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__5__0_chanx_left_out[0:228]),
		.ccff_tail(sb_3__5__0_ccff_tail));

	sb_3__5_ sb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__4_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_4_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_4_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__5__4_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__5_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_3__5__1_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_4_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__4_ccff_tail),
		.chany_top_out(sb_3__5__1_chany_top_out[0:228]),
		.chanx_right_out(sb_3__5__1_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__5__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__5__1_chanx_left_out[0:228]),
		.ccff_tail(sb_3__5__1_ccff_tail));

	sb_3__5_ sb_9__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__3__7_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_7_right_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_oack_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_7_right_width_0_height_0_subtile_0__pin_olck_1_1_),
		.chanx_right_in(cbx_1__5__6_chanx_left_out[0:228]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_16_),
		.chany_bottom_in(cby_1__5__8_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_3__5__2_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_7_bottom_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(cbx_1__5__6_ccff_tail),
		.chany_top_out(sb_3__5__2_chany_top_out[0:228]),
		.chanx_right_out(sb_3__5__2_chanx_right_out[0:228]),
		.chany_bottom_out(sb_3__5__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_3__5__2_chanx_left_out[0:228]),
		.ccff_tail(sb_3__5__2_ccff_tail));

	sb_22__0_ sb_22__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__0_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__21_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(cbx_1__0__20_ccff_tail),
		.chany_top_out(sb_22__0__0_chany_top_out[0:228]),
		.chanx_left_out(sb_22__0__0_chanx_left_out[0:228]),
		.ccff_tail(sb_22__0__0_ccff_tail));

	sb_22__1_ sb_22__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__1_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__0_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_21_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__384_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__0_ccff_tail),
		.chany_top_out(sb_22__1__0_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__0_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__0_ccff_tail));

	sb_22__1_ sb_22__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__2_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__1_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_20_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__385_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__351_ccff_tail),
		.chany_top_out(sb_22__1__1_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__1_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__1_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__1_ccff_tail));

	sb_22__1_ sb_22__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__3_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__2_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__386_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__2_ccff_tail),
		.chany_top_out(sb_22__1__2_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__2_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__2_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__2_ccff_tail));

	sb_22__1_ sb_22__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__5_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__4_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__387_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__353_ccff_tail),
		.chany_top_out(sb_22__1__3_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__3_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__3_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__3_ccff_tail));

	sb_22__1_ sb_22__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__6_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__5_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__388_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__5_ccff_tail),
		.chany_top_out(sb_22__1__4_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__4_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__4_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__4_ccff_tail));

	sb_22__1_ sb_22__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__7_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__6_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__389_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__355_ccff_tail),
		.chany_top_out(sb_22__1__5_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__5_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__5_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__5_ccff_tail));

	sb_22__1_ sb_22__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__8_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__7_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__390_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__7_ccff_tail),
		.chany_top_out(sb_22__1__6_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__6_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__6_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__6_ccff_tail));

	sb_22__1_ sb_22__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__9_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__8_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__391_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__357_ccff_tail),
		.chany_top_out(sb_22__1__7_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__7_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__7_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__7_ccff_tail));

	sb_22__1_ sb_22__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__10_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__9_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__392_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__9_ccff_tail),
		.chany_top_out(sb_22__1__8_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__8_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__8_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__8_ccff_tail));

	sb_22__1_ sb_22__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__11_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__10_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__393_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__359_ccff_tail),
		.chany_top_out(sb_22__1__9_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__9_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__9_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__9_ccff_tail));

	sb_22__1_ sb_22__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__12_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__11_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__394_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__11_ccff_tail),
		.chany_top_out(sb_22__1__10_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__10_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__10_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__10_ccff_tail));

	sb_22__1_ sb_22__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__13_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__12_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__395_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__361_ccff_tail),
		.chany_top_out(sb_22__1__11_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__11_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__11_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__11_ccff_tail));

	sb_22__1_ sb_22__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__14_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__13_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__396_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__13_ccff_tail),
		.chany_top_out(sb_22__1__12_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__12_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__12_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__12_ccff_tail));

	sb_22__1_ sb_22__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__15_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__14_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__397_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__363_ccff_tail),
		.chany_top_out(sb_22__1__13_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__13_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__13_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__13_ccff_tail));

	sb_22__1_ sb_22__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__16_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__15_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__398_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__15_ccff_tail),
		.chany_top_out(sb_22__1__14_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__14_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__14_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__14_ccff_tail));

	sb_22__1_ sb_22__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__17_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__16_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__399_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__365_ccff_tail),
		.chany_top_out(sb_22__1__15_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__15_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__15_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__15_ccff_tail));

	sb_22__1_ sb_22__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__18_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__17_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__400_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__17_ccff_tail),
		.chany_top_out(sb_22__1__16_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__16_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__16_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__16_ccff_tail));

	sb_22__1_ sb_22__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__19_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__18_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__401_chanx_right_out[0:228]),
		.ccff_head(sb_1__1__367_ccff_tail),
		.chany_top_out(sb_22__1__17_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__17_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__17_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__17_ccff_tail));

	sb_22__1_ sb_22__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__20_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__19_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__1__402_chanx_right_out[0:228]),
		.ccff_head(cby_22__1__19_ccff_tail),
		.chany_top_out(sb_22__1__18_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__1__18_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__1__18_chanx_left_out[0:228]),
		.ccff_tail(sb_22__1__18_ccff_tail));

	sb_22__4_ sb_22__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__5__0_chany_bottom_out[0:228]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__1__3_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__4__21_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_22__4__0_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__4__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__4__0_chanx_left_out[0:228]),
		.ccff_tail(sb_22__4__0_ccff_tail));

	sb_22__5_ sb_22__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_22__1__4_chany_bottom_out[0:228]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_22__5__0_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.chanx_left_in(cbx_1__5__18_chanx_right_out[0:228]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_16_),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_22__5__0_chany_top_out[0:228]),
		.chany_bottom_out(sb_22__5__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__5__0_chanx_left_out[0:228]),
		.ccff_tail(sb_22__5__0_ccff_tail));

	sb_22__22_ sb_22__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_22__1__20_chany_top_out[0:228]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__22__21_chanx_right_out[0:228]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_21_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_22__22__0_chany_bottom_out[0:228]),
		.chanx_left_out(sb_22__22__0_chanx_left_out[0:228]),
		.ccff_tail(sb_22__22__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__5_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__6_ccff_tail),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__6_ccff_tail));

	cbx_1__0_ cbx_8__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__7_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__7_ccff_tail),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__7_ccff_tail));

	cbx_1__0_ cbx_9__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__8_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__8_ccff_tail),
		.chanx_left_out(cbx_1__0__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__8_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__8_ccff_tail));

	cbx_1__0_ cbx_10__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__9_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__9_ccff_tail),
		.chanx_left_out(cbx_1__0__9_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__9_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__9_ccff_tail));

	cbx_1__0_ cbx_11__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__10_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__10_ccff_tail),
		.chanx_left_out(cbx_1__0__10_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__10_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__10_ccff_tail));

	cbx_1__0_ cbx_12__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__11_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__11_ccff_tail),
		.chanx_left_out(cbx_1__0__11_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__11_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__11_ccff_tail));

	cbx_1__0_ cbx_13__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__12_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__12_ccff_tail),
		.chanx_left_out(cbx_1__0__12_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__12_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__12_ccff_tail));

	cbx_1__0_ cbx_14__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__13_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__13_ccff_tail),
		.chanx_left_out(cbx_1__0__13_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__13_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__13_ccff_tail));

	cbx_1__0_ cbx_15__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__14_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__14_ccff_tail),
		.chanx_left_out(cbx_1__0__14_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__14_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__14_ccff_tail));

	cbx_1__0_ cbx_16__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__15_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__15_ccff_tail),
		.chanx_left_out(cbx_1__0__15_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__15_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__15_ccff_tail));

	cbx_1__0_ cbx_17__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__15_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__16_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__16_ccff_tail),
		.chanx_left_out(cbx_1__0__16_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__16_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__16_ccff_tail));

	cbx_1__0_ cbx_18__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__16_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__17_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__17_ccff_tail),
		.chanx_left_out(cbx_1__0__17_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__17_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__17_ccff_tail));

	cbx_1__0_ cbx_19__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__17_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__18_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__18_ccff_tail),
		.chanx_left_out(cbx_1__0__18_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__18_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__18_ccff_tail));

	cbx_1__0_ cbx_20__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__18_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__19_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__19_ccff_tail),
		.chanx_left_out(cbx_1__0__19_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__19_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__19_ccff_tail));

	cbx_1__0_ cbx_21__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__19_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__0__20_chanx_left_out[0:228]),
		.ccff_head(sb_1__0__20_ccff_tail),
		.chanx_left_out(cbx_1__0__20_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__20_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__20_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__20_ccff_tail));

	cbx_1__0_ cbx_22__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__20_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__0__0_chanx_left_out[0:228]),
		.ccff_head(sb_22__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__21_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__0__21_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__21_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__21_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__2_ (
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__3_ (
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__6_ (
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__7_ (
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__8_ (
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__9_ (
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__10_ (
		.chanx_left_in(sb_0__1__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__11_ (
		.chanx_left_in(sb_0__1__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__12_ (
		.chanx_left_in(sb_0__1__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__13_ (
		.chanx_left_in(sb_0__1__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__14_ (
		.chanx_left_in(sb_0__1__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__15_ (
		.chanx_left_in(sb_0__1__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__16_ (
		.chanx_left_in(sb_0__1__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__17_ (
		.chanx_left_in(sb_0__1__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__18_ (
		.chanx_left_in(sb_0__1__15_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__19_ (
		.chanx_left_in(sb_0__1__16_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__20_ (
		.chanx_left_in(sb_0__1__17_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:228]));

	cbx_1__1_ cbx_1__21_ (
		.chanx_left_in(sb_0__1__18_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__1_ (
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__2_ (
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__0_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__20_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__20_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__3_ (
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__0_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__21_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__21_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__6_ (
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__1_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__22_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__22_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__7_ (
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__23_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__23_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__8_ (
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__1_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__24_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__24_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__9_ (
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__2_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__25_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__25_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__10_ (
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__26_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__26_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__11_ (
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__27_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__27_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__12_ (
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__28_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__28_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__13_ (
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__29_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__29_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__14_ (
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__30_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__30_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__15_ (
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__31_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__31_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__16_ (
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__32_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__32_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__17_ (
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__33_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__33_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__18_ (
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__34_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__34_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__19_ (
		.chanx_left_in(sb_1__1__16_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__35_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__35_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__20_ (
		.chanx_left_in(sb_1__1__17_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__36_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__36_chanx_right_out[0:228]));

	cbx_1__1_ cbx_2__21_ (
		.chanx_left_in(sb_1__1__18_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__37_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__37_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__1_ (
		.chanx_left_in(sb_1__1__19_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__38_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__38_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__7_ (
		.chanx_left_in(sb_1__1__20_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__39_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__39_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__10_ (
		.chanx_left_in(sb_1__1__21_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__40_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__40_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__11_ (
		.chanx_left_in(sb_1__1__22_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__41_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__41_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__12_ (
		.chanx_left_in(sb_1__1__23_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__42_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__42_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__13_ (
		.chanx_left_in(sb_1__1__24_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__43_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__43_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__14_ (
		.chanx_left_in(sb_1__1__25_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__44_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__44_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__15_ (
		.chanx_left_in(sb_1__1__26_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__45_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__45_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__16_ (
		.chanx_left_in(sb_1__1__27_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__46_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__46_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__17_ (
		.chanx_left_in(sb_1__1__28_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__47_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__47_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__18_ (
		.chanx_left_in(sb_1__1__29_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__48_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__48_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__19_ (
		.chanx_left_in(sb_1__1__30_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__49_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__49_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__20_ (
		.chanx_left_in(sb_1__1__31_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__50_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__50_chanx_right_out[0:228]));

	cbx_1__1_ cbx_3__21_ (
		.chanx_left_in(sb_1__1__32_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__51_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__51_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__1_ (
		.chanx_left_in(sb_1__1__33_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__52_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__52_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__2_ (
		.chanx_left_in(sb_3__2__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__53_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__53_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__3_ (
		.chanx_left_in(sb_3__3__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__49_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__54_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__54_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__6_ (
		.chanx_left_in(sb_3__3__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__50_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__55_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__55_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__7_ (
		.chanx_left_in(sb_1__1__34_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__51_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__56_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__56_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__8_ (
		.chanx_left_in(sb_3__2__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__52_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__57_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__57_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__9_ (
		.chanx_left_in(sb_3__3__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__53_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__58_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__58_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__10_ (
		.chanx_left_in(sb_1__1__35_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__54_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__59_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__59_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__11_ (
		.chanx_left_in(sb_1__1__36_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__55_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__60_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__60_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__12_ (
		.chanx_left_in(sb_1__1__37_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__56_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__61_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__61_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__13_ (
		.chanx_left_in(sb_1__1__38_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__57_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__62_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__62_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__14_ (
		.chanx_left_in(sb_1__1__39_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__58_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__63_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__63_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__15_ (
		.chanx_left_in(sb_1__1__40_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__59_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__64_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__64_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__16_ (
		.chanx_left_in(sb_1__1__41_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__60_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__65_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__65_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__17_ (
		.chanx_left_in(sb_1__1__42_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__61_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__66_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__66_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__18_ (
		.chanx_left_in(sb_1__1__43_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__62_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__67_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__67_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__19_ (
		.chanx_left_in(sb_1__1__44_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__63_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__68_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__68_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__20_ (
		.chanx_left_in(sb_1__1__45_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__64_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__69_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__69_chanx_right_out[0:228]));

	cbx_1__1_ cbx_4__21_ (
		.chanx_left_in(sb_1__1__46_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__65_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__70_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__70_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__1_ (
		.chanx_left_in(sb_1__1__47_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__66_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__71_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__71_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__2_ (
		.chanx_left_in(sb_1__1__48_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__2_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__72_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__72_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__3_ (
		.chanx_left_in(sb_1__1__49_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__3_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__73_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__73_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__6_ (
		.chanx_left_in(sb_1__1__50_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__4_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__74_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__74_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__7_ (
		.chanx_left_in(sb_1__1__51_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__67_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__75_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__75_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__8_ (
		.chanx_left_in(sb_1__1__52_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__3_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__76_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__76_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__9_ (
		.chanx_left_in(sb_1__1__53_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__5_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__77_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__77_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__10_ (
		.chanx_left_in(sb_1__1__54_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__68_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__78_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__78_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__11_ (
		.chanx_left_in(sb_1__1__55_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__69_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__79_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__79_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__12_ (
		.chanx_left_in(sb_1__1__56_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__70_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__80_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__80_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__13_ (
		.chanx_left_in(sb_1__1__57_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__71_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__81_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__81_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__14_ (
		.chanx_left_in(sb_1__1__58_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__72_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__82_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__82_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__15_ (
		.chanx_left_in(sb_1__1__59_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__73_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__83_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__83_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__16_ (
		.chanx_left_in(sb_1__1__60_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__74_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__84_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__84_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__17_ (
		.chanx_left_in(sb_1__1__61_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__75_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__85_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__85_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__18_ (
		.chanx_left_in(sb_1__1__62_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__76_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__86_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__86_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__19_ (
		.chanx_left_in(sb_1__1__63_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__77_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__87_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__87_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__20_ (
		.chanx_left_in(sb_1__1__64_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__78_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__88_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__88_chanx_right_out[0:228]));

	cbx_1__1_ cbx_5__21_ (
		.chanx_left_in(sb_1__1__65_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__79_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__89_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__89_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__1_ (
		.chanx_left_in(sb_1__1__66_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__80_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__90_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__90_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__7_ (
		.chanx_left_in(sb_1__1__67_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__81_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__91_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__91_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__10_ (
		.chanx_left_in(sb_1__1__68_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__82_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__92_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__92_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__11_ (
		.chanx_left_in(sb_1__1__69_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__83_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__93_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__93_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__12_ (
		.chanx_left_in(sb_1__1__70_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__84_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__94_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__94_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__13_ (
		.chanx_left_in(sb_1__1__71_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__85_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__95_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__95_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__14_ (
		.chanx_left_in(sb_1__1__72_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__86_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__96_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__96_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__15_ (
		.chanx_left_in(sb_1__1__73_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__87_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__97_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__97_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__16_ (
		.chanx_left_in(sb_1__1__74_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__88_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__98_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__98_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__17_ (
		.chanx_left_in(sb_1__1__75_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__89_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__99_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__99_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__18_ (
		.chanx_left_in(sb_1__1__76_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__90_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__100_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__100_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__19_ (
		.chanx_left_in(sb_1__1__77_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__91_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__101_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__101_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__20_ (
		.chanx_left_in(sb_1__1__78_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__92_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__102_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__102_chanx_right_out[0:228]));

	cbx_1__1_ cbx_6__21_ (
		.chanx_left_in(sb_1__1__79_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__93_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__103_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__103_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__1_ (
		.chanx_left_in(sb_1__1__80_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__94_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__104_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__104_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__2_ (
		.chanx_left_in(sb_3__2__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__95_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__105_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__105_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__3_ (
		.chanx_left_in(sb_3__3__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__96_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__106_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__106_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__6_ (
		.chanx_left_in(sb_3__3__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__97_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__107_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__107_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__7_ (
		.chanx_left_in(sb_1__1__81_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__98_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__108_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__108_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__8_ (
		.chanx_left_in(sb_3__2__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__99_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__109_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__109_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__9_ (
		.chanx_left_in(sb_3__3__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__100_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__110_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__110_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__10_ (
		.chanx_left_in(sb_1__1__82_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__101_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__111_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__111_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__11_ (
		.chanx_left_in(sb_1__1__83_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__102_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__112_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__112_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__12_ (
		.chanx_left_in(sb_1__1__84_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__103_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__113_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__113_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__13_ (
		.chanx_left_in(sb_1__1__85_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__104_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__114_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__114_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__14_ (
		.chanx_left_in(sb_1__1__86_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__105_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__115_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__115_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__15_ (
		.chanx_left_in(sb_1__1__87_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__106_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__116_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__116_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__16_ (
		.chanx_left_in(sb_1__1__88_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__107_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__117_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__117_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__17_ (
		.chanx_left_in(sb_1__1__89_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__108_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__118_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__118_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__18_ (
		.chanx_left_in(sb_1__1__90_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__109_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__119_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__119_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__19_ (
		.chanx_left_in(sb_1__1__91_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__110_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__120_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__120_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__20_ (
		.chanx_left_in(sb_1__1__92_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__111_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__121_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__121_chanx_right_out[0:228]));

	cbx_1__1_ cbx_7__21_ (
		.chanx_left_in(sb_1__1__93_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__112_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__122_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__122_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__1_ (
		.chanx_left_in(sb_1__1__94_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__113_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__123_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__123_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__2_ (
		.chanx_left_in(sb_1__1__95_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__4_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__124_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__124_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__3_ (
		.chanx_left_in(sb_1__1__96_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__6_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__125_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__125_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__6_ (
		.chanx_left_in(sb_1__1__97_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__7_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__126_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__126_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__7_ (
		.chanx_left_in(sb_1__1__98_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__114_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__127_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__127_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__8_ (
		.chanx_left_in(sb_1__1__99_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__2__5_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__128_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__128_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__9_ (
		.chanx_left_in(sb_1__1__100_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__3__8_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__129_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__129_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__10_ (
		.chanx_left_in(sb_1__1__101_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__115_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__130_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__130_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__11_ (
		.chanx_left_in(sb_1__1__102_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__116_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__131_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__131_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__12_ (
		.chanx_left_in(sb_1__1__103_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__117_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__132_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__132_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__13_ (
		.chanx_left_in(sb_1__1__104_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__118_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__133_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__133_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__14_ (
		.chanx_left_in(sb_1__1__105_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__119_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__134_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__134_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__15_ (
		.chanx_left_in(sb_1__1__106_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__120_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__135_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__135_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__16_ (
		.chanx_left_in(sb_1__1__107_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__121_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__136_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__136_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__17_ (
		.chanx_left_in(sb_1__1__108_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__122_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__137_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__137_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__18_ (
		.chanx_left_in(sb_1__1__109_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__123_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__138_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__138_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__19_ (
		.chanx_left_in(sb_1__1__110_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__124_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__139_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__139_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__20_ (
		.chanx_left_in(sb_1__1__111_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__125_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__140_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__140_chanx_right_out[0:228]));

	cbx_1__1_ cbx_8__21_ (
		.chanx_left_in(sb_1__1__112_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__126_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__141_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__141_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__1_ (
		.chanx_left_in(sb_1__1__113_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__127_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__142_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__142_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__7_ (
		.chanx_left_in(sb_1__1__114_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__128_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__143_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__143_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__10_ (
		.chanx_left_in(sb_1__1__115_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__129_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__144_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__144_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__11_ (
		.chanx_left_in(sb_1__1__116_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__130_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__145_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__145_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__12_ (
		.chanx_left_in(sb_1__1__117_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__131_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__146_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__146_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__13_ (
		.chanx_left_in(sb_1__1__118_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__132_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__147_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__147_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__14_ (
		.chanx_left_in(sb_1__1__119_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__133_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__148_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__148_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__15_ (
		.chanx_left_in(sb_1__1__120_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__134_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__149_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__149_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__16_ (
		.chanx_left_in(sb_1__1__121_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__135_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__150_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__150_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__17_ (
		.chanx_left_in(sb_1__1__122_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__136_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__151_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__151_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__18_ (
		.chanx_left_in(sb_1__1__123_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__137_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__152_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__152_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__19_ (
		.chanx_left_in(sb_1__1__124_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__138_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__153_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__153_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__20_ (
		.chanx_left_in(sb_1__1__125_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__139_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__154_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__154_chanx_right_out[0:228]));

	cbx_1__1_ cbx_9__21_ (
		.chanx_left_in(sb_1__1__126_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__140_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__155_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__155_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__1_ (
		.chanx_left_in(sb_1__1__127_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__141_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__156_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__156_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__2_ (
		.chanx_left_in(sb_3__2__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__142_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__157_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__157_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__3_ (
		.chanx_left_in(sb_3__3__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__143_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__158_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__158_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__6_ (
		.chanx_left_in(sb_3__3__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__144_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__159_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__159_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__7_ (
		.chanx_left_in(sb_1__1__128_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__145_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__160_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__160_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__8_ (
		.chanx_left_in(sb_3__2__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__146_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__161_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__161_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__9_ (
		.chanx_left_in(sb_3__3__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__147_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__162_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__162_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__10_ (
		.chanx_left_in(sb_1__1__129_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__148_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__163_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__163_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__11_ (
		.chanx_left_in(sb_1__1__130_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__149_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__164_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__164_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__12_ (
		.chanx_left_in(sb_1__1__131_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__150_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__165_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__165_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__13_ (
		.chanx_left_in(sb_1__1__132_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__151_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__166_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__166_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__14_ (
		.chanx_left_in(sb_1__1__133_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__152_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__167_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__167_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__15_ (
		.chanx_left_in(sb_1__1__134_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__153_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__168_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__168_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__16_ (
		.chanx_left_in(sb_1__1__135_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__154_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__169_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__169_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__17_ (
		.chanx_left_in(sb_1__1__136_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__155_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__170_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__170_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__18_ (
		.chanx_left_in(sb_1__1__137_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__156_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__171_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__171_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__19_ (
		.chanx_left_in(sb_1__1__138_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__157_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__172_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__172_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__20_ (
		.chanx_left_in(sb_1__1__139_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__158_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__173_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__173_chanx_right_out[0:228]));

	cbx_1__1_ cbx_10__21_ (
		.chanx_left_in(sb_1__1__140_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__159_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__174_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__174_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__1_ (
		.chanx_left_in(sb_1__1__141_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__160_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__175_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__175_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__2_ (
		.chanx_left_in(sb_1__1__142_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__161_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__176_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__176_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__3_ (
		.chanx_left_in(sb_1__1__143_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__162_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__177_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__177_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__6_ (
		.chanx_left_in(sb_1__1__144_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__163_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__178_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__178_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__7_ (
		.chanx_left_in(sb_1__1__145_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__164_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__179_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__179_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__8_ (
		.chanx_left_in(sb_1__1__146_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__165_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__180_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__180_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__9_ (
		.chanx_left_in(sb_1__1__147_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__166_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__181_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__181_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__10_ (
		.chanx_left_in(sb_1__1__148_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__167_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__182_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__182_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__11_ (
		.chanx_left_in(sb_1__1__149_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__168_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__183_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__183_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__12_ (
		.chanx_left_in(sb_1__1__150_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__169_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__184_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__184_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__13_ (
		.chanx_left_in(sb_1__1__151_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__170_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__185_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__185_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__14_ (
		.chanx_left_in(sb_1__1__152_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__171_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__186_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__186_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__15_ (
		.chanx_left_in(sb_1__1__153_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__172_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__187_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__187_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__16_ (
		.chanx_left_in(sb_1__1__154_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__173_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__188_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__188_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__17_ (
		.chanx_left_in(sb_1__1__155_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__174_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__189_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__189_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__18_ (
		.chanx_left_in(sb_1__1__156_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__175_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__190_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__190_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__19_ (
		.chanx_left_in(sb_1__1__157_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__176_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__191_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__191_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__20_ (
		.chanx_left_in(sb_1__1__158_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__177_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__192_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__192_chanx_right_out[0:228]));

	cbx_1__1_ cbx_11__21_ (
		.chanx_left_in(sb_1__1__159_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__178_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__193_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__193_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__1_ (
		.chanx_left_in(sb_1__1__160_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__179_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__194_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__194_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__2_ (
		.chanx_left_in(sb_1__1__161_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__180_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__195_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__195_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__3_ (
		.chanx_left_in(sb_1__1__162_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__181_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__196_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__196_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__6_ (
		.chanx_left_in(sb_1__1__163_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__182_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__197_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__197_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__7_ (
		.chanx_left_in(sb_1__1__164_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__183_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__198_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__198_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__8_ (
		.chanx_left_in(sb_1__1__165_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__184_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__199_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__199_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__9_ (
		.chanx_left_in(sb_1__1__166_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__185_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__200_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__200_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__10_ (
		.chanx_left_in(sb_1__1__167_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__186_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__201_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__201_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__11_ (
		.chanx_left_in(sb_1__1__168_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__187_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__202_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__202_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__12_ (
		.chanx_left_in(sb_1__1__169_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__188_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__203_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__203_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__13_ (
		.chanx_left_in(sb_1__1__170_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__189_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__204_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__204_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__14_ (
		.chanx_left_in(sb_1__1__171_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__190_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__205_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__205_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__15_ (
		.chanx_left_in(sb_1__1__172_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__191_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__206_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__206_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__16_ (
		.chanx_left_in(sb_1__1__173_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__192_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__207_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__207_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__17_ (
		.chanx_left_in(sb_1__1__174_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__193_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__208_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__208_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__18_ (
		.chanx_left_in(sb_1__1__175_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__194_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__209_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__209_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__19_ (
		.chanx_left_in(sb_1__1__176_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__195_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__210_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__210_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__20_ (
		.chanx_left_in(sb_1__1__177_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__196_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__211_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__211_chanx_right_out[0:228]));

	cbx_1__1_ cbx_12__21_ (
		.chanx_left_in(sb_1__1__178_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__197_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__212_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__212_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__1_ (
		.chanx_left_in(sb_1__1__179_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__198_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__213_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__213_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__2_ (
		.chanx_left_in(sb_1__1__180_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__199_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__214_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__214_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__3_ (
		.chanx_left_in(sb_1__1__181_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__200_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__215_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__215_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__6_ (
		.chanx_left_in(sb_1__1__182_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__201_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__216_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__216_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__7_ (
		.chanx_left_in(sb_1__1__183_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__202_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__217_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__217_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__8_ (
		.chanx_left_in(sb_1__1__184_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__203_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__218_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__218_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__9_ (
		.chanx_left_in(sb_1__1__185_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__204_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__219_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__219_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__10_ (
		.chanx_left_in(sb_1__1__186_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__205_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__220_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__220_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__11_ (
		.chanx_left_in(sb_1__1__187_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__206_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__221_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__221_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__12_ (
		.chanx_left_in(sb_1__1__188_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__207_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__222_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__222_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__13_ (
		.chanx_left_in(sb_1__1__189_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__208_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__223_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__223_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__14_ (
		.chanx_left_in(sb_1__1__190_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__209_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__224_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__224_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__15_ (
		.chanx_left_in(sb_1__1__191_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__210_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__225_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__225_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__16_ (
		.chanx_left_in(sb_1__1__192_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__211_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__226_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__226_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__17_ (
		.chanx_left_in(sb_1__1__193_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__212_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__227_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__227_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__18_ (
		.chanx_left_in(sb_1__1__194_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__213_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__228_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__228_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__19_ (
		.chanx_left_in(sb_1__1__195_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__214_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__229_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__229_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__20_ (
		.chanx_left_in(sb_1__1__196_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__215_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__230_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__230_chanx_right_out[0:228]));

	cbx_1__1_ cbx_13__21_ (
		.chanx_left_in(sb_1__1__197_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__216_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__231_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__231_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__1_ (
		.chanx_left_in(sb_1__1__198_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__217_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__232_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__232_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__2_ (
		.chanx_left_in(sb_1__1__199_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__218_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__233_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__233_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__3_ (
		.chanx_left_in(sb_1__1__200_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__219_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__234_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__234_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__6_ (
		.chanx_left_in(sb_1__1__201_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__220_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__235_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__235_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__7_ (
		.chanx_left_in(sb_1__1__202_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__221_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__236_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__236_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__8_ (
		.chanx_left_in(sb_1__1__203_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__222_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__237_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__237_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__9_ (
		.chanx_left_in(sb_1__1__204_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__223_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__238_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__238_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__10_ (
		.chanx_left_in(sb_1__1__205_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__224_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__239_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__239_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__11_ (
		.chanx_left_in(sb_1__1__206_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__225_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__240_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__240_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__12_ (
		.chanx_left_in(sb_1__1__207_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__226_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__241_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__241_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__13_ (
		.chanx_left_in(sb_1__1__208_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__227_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__242_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__242_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__14_ (
		.chanx_left_in(sb_1__1__209_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__228_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__243_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__243_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__15_ (
		.chanx_left_in(sb_1__1__210_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__229_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__244_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__244_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__16_ (
		.chanx_left_in(sb_1__1__211_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__230_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__245_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__245_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__17_ (
		.chanx_left_in(sb_1__1__212_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__231_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__246_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__246_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__18_ (
		.chanx_left_in(sb_1__1__213_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__232_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__247_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__247_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__19_ (
		.chanx_left_in(sb_1__1__214_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__233_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__248_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__248_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__20_ (
		.chanx_left_in(sb_1__1__215_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__234_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__249_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__249_chanx_right_out[0:228]));

	cbx_1__1_ cbx_14__21_ (
		.chanx_left_in(sb_1__1__216_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__235_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__250_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__250_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__1_ (
		.chanx_left_in(sb_1__1__217_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__236_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__251_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__251_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__2_ (
		.chanx_left_in(sb_1__1__218_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__237_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__252_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__252_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__3_ (
		.chanx_left_in(sb_1__1__219_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__238_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__253_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__253_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__6_ (
		.chanx_left_in(sb_1__1__220_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__239_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__254_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__254_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__7_ (
		.chanx_left_in(sb_1__1__221_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__240_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__255_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__255_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__8_ (
		.chanx_left_in(sb_1__1__222_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__241_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__256_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__256_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__9_ (
		.chanx_left_in(sb_1__1__223_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__242_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__257_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__257_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__10_ (
		.chanx_left_in(sb_1__1__224_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__243_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__258_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__258_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__11_ (
		.chanx_left_in(sb_1__1__225_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__244_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__259_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__259_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__12_ (
		.chanx_left_in(sb_1__1__226_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__245_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__260_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__260_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__13_ (
		.chanx_left_in(sb_1__1__227_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__246_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__261_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__261_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__14_ (
		.chanx_left_in(sb_1__1__228_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__247_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__262_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__262_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__15_ (
		.chanx_left_in(sb_1__1__229_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__248_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__263_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__263_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__16_ (
		.chanx_left_in(sb_1__1__230_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__249_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__264_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__264_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__17_ (
		.chanx_left_in(sb_1__1__231_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__250_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__265_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__265_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__18_ (
		.chanx_left_in(sb_1__1__232_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__251_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__266_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__266_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__19_ (
		.chanx_left_in(sb_1__1__233_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__252_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__267_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__267_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__20_ (
		.chanx_left_in(sb_1__1__234_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__253_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__268_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__268_chanx_right_out[0:228]));

	cbx_1__1_ cbx_15__21_ (
		.chanx_left_in(sb_1__1__235_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__254_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__269_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__269_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__1_ (
		.chanx_left_in(sb_1__1__236_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__255_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__270_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__270_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__2_ (
		.chanx_left_in(sb_1__1__237_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__256_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__271_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__271_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__3_ (
		.chanx_left_in(sb_1__1__238_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__257_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__272_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__272_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__6_ (
		.chanx_left_in(sb_1__1__239_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__258_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__273_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__273_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__7_ (
		.chanx_left_in(sb_1__1__240_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__259_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__274_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__274_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__8_ (
		.chanx_left_in(sb_1__1__241_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__260_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__275_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__275_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__9_ (
		.chanx_left_in(sb_1__1__242_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__261_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__276_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__276_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__10_ (
		.chanx_left_in(sb_1__1__243_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__262_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__277_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__277_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__11_ (
		.chanx_left_in(sb_1__1__244_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__263_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__278_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__278_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__12_ (
		.chanx_left_in(sb_1__1__245_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__264_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__279_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__279_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__13_ (
		.chanx_left_in(sb_1__1__246_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__265_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__280_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__280_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__14_ (
		.chanx_left_in(sb_1__1__247_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__266_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__281_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__281_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__15_ (
		.chanx_left_in(sb_1__1__248_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__267_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__282_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__282_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__16_ (
		.chanx_left_in(sb_1__1__249_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__268_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__283_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__283_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__17_ (
		.chanx_left_in(sb_1__1__250_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__269_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__284_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__284_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__18_ (
		.chanx_left_in(sb_1__1__251_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__270_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__285_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__285_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__19_ (
		.chanx_left_in(sb_1__1__252_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__271_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__286_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__286_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__20_ (
		.chanx_left_in(sb_1__1__253_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__272_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__287_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__287_chanx_right_out[0:228]));

	cbx_1__1_ cbx_16__21_ (
		.chanx_left_in(sb_1__1__254_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__273_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__288_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__288_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__1_ (
		.chanx_left_in(sb_1__1__255_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__274_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__289_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__289_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__2_ (
		.chanx_left_in(sb_1__1__256_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__275_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__290_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__290_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__3_ (
		.chanx_left_in(sb_1__1__257_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__276_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__291_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__291_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__6_ (
		.chanx_left_in(sb_1__1__258_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__277_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__292_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__292_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__7_ (
		.chanx_left_in(sb_1__1__259_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__278_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__293_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__293_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__8_ (
		.chanx_left_in(sb_1__1__260_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__279_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__294_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__294_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__9_ (
		.chanx_left_in(sb_1__1__261_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__280_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__295_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__295_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__10_ (
		.chanx_left_in(sb_1__1__262_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__281_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__296_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__296_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__11_ (
		.chanx_left_in(sb_1__1__263_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__282_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__297_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__297_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__12_ (
		.chanx_left_in(sb_1__1__264_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__283_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__298_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__298_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__13_ (
		.chanx_left_in(sb_1__1__265_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__284_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__299_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__299_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__14_ (
		.chanx_left_in(sb_1__1__266_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__285_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__300_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__300_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__15_ (
		.chanx_left_in(sb_1__1__267_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__286_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__301_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__301_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__16_ (
		.chanx_left_in(sb_1__1__268_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__287_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__302_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__302_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__17_ (
		.chanx_left_in(sb_1__1__269_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__288_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__303_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__303_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__18_ (
		.chanx_left_in(sb_1__1__270_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__289_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__304_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__304_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__19_ (
		.chanx_left_in(sb_1__1__271_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__290_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__305_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__305_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__20_ (
		.chanx_left_in(sb_1__1__272_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__291_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__306_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__306_chanx_right_out[0:228]));

	cbx_1__1_ cbx_17__21_ (
		.chanx_left_in(sb_1__1__273_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__292_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__307_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__307_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__1_ (
		.chanx_left_in(sb_1__1__274_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__293_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__308_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__308_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__2_ (
		.chanx_left_in(sb_1__1__275_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__294_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__309_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__309_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__3_ (
		.chanx_left_in(sb_1__1__276_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__295_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__310_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__310_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__6_ (
		.chanx_left_in(sb_1__1__277_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__296_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__311_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__311_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__7_ (
		.chanx_left_in(sb_1__1__278_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__297_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__312_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__312_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__8_ (
		.chanx_left_in(sb_1__1__279_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__298_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__313_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__313_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__9_ (
		.chanx_left_in(sb_1__1__280_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__299_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__314_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__314_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__10_ (
		.chanx_left_in(sb_1__1__281_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__300_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__315_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__315_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__11_ (
		.chanx_left_in(sb_1__1__282_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__301_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__316_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__316_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__12_ (
		.chanx_left_in(sb_1__1__283_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__302_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__317_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__317_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__13_ (
		.chanx_left_in(sb_1__1__284_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__303_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__318_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__318_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__14_ (
		.chanx_left_in(sb_1__1__285_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__304_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__319_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__319_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__15_ (
		.chanx_left_in(sb_1__1__286_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__305_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__320_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__320_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__16_ (
		.chanx_left_in(sb_1__1__287_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__306_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__321_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__321_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__17_ (
		.chanx_left_in(sb_1__1__288_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__307_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__322_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__322_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__18_ (
		.chanx_left_in(sb_1__1__289_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__308_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__323_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__323_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__19_ (
		.chanx_left_in(sb_1__1__290_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__309_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__324_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__324_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__20_ (
		.chanx_left_in(sb_1__1__291_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__310_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__325_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__325_chanx_right_out[0:228]));

	cbx_1__1_ cbx_18__21_ (
		.chanx_left_in(sb_1__1__292_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__311_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__326_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__326_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__1_ (
		.chanx_left_in(sb_1__1__293_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__312_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__327_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__327_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__2_ (
		.chanx_left_in(sb_1__1__294_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__313_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__328_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__328_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__3_ (
		.chanx_left_in(sb_1__1__295_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__314_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__329_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__329_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__6_ (
		.chanx_left_in(sb_1__1__296_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__315_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__330_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__330_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__7_ (
		.chanx_left_in(sb_1__1__297_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__316_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__331_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__331_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__8_ (
		.chanx_left_in(sb_1__1__298_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__317_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__332_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__332_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__9_ (
		.chanx_left_in(sb_1__1__299_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__318_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__333_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__333_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__10_ (
		.chanx_left_in(sb_1__1__300_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__319_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__334_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__334_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__11_ (
		.chanx_left_in(sb_1__1__301_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__320_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__335_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__335_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__12_ (
		.chanx_left_in(sb_1__1__302_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__321_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__336_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__336_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__13_ (
		.chanx_left_in(sb_1__1__303_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__322_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__337_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__337_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__14_ (
		.chanx_left_in(sb_1__1__304_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__323_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__338_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__338_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__15_ (
		.chanx_left_in(sb_1__1__305_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__324_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__339_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__339_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__16_ (
		.chanx_left_in(sb_1__1__306_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__325_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__340_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__340_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__17_ (
		.chanx_left_in(sb_1__1__307_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__326_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__341_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__341_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__18_ (
		.chanx_left_in(sb_1__1__308_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__327_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__342_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__342_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__19_ (
		.chanx_left_in(sb_1__1__309_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__328_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__343_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__343_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__20_ (
		.chanx_left_in(sb_1__1__310_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__329_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__344_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__344_chanx_right_out[0:228]));

	cbx_1__1_ cbx_19__21_ (
		.chanx_left_in(sb_1__1__311_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__330_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__345_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__345_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__1_ (
		.chanx_left_in(sb_1__1__312_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__331_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__346_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__346_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__2_ (
		.chanx_left_in(sb_1__1__313_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__332_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__347_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__347_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__3_ (
		.chanx_left_in(sb_1__1__314_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__333_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__348_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__348_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__6_ (
		.chanx_left_in(sb_1__1__315_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__334_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__349_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__349_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__7_ (
		.chanx_left_in(sb_1__1__316_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__335_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__350_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__350_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__8_ (
		.chanx_left_in(sb_1__1__317_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__336_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__351_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__351_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__9_ (
		.chanx_left_in(sb_1__1__318_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__337_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__352_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__352_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__10_ (
		.chanx_left_in(sb_1__1__319_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__338_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__353_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__353_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__11_ (
		.chanx_left_in(sb_1__1__320_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__339_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__354_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__354_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__12_ (
		.chanx_left_in(sb_1__1__321_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__340_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__355_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__355_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__13_ (
		.chanx_left_in(sb_1__1__322_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__341_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__356_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__356_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__14_ (
		.chanx_left_in(sb_1__1__323_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__342_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__357_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__357_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__15_ (
		.chanx_left_in(sb_1__1__324_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__343_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__358_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__358_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__16_ (
		.chanx_left_in(sb_1__1__325_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__344_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__359_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__359_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__17_ (
		.chanx_left_in(sb_1__1__326_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__345_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__360_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__360_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__18_ (
		.chanx_left_in(sb_1__1__327_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__346_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__361_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__361_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__19_ (
		.chanx_left_in(sb_1__1__328_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__347_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__362_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__362_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__20_ (
		.chanx_left_in(sb_1__1__329_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__348_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__363_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__363_chanx_right_out[0:228]));

	cbx_1__1_ cbx_20__21_ (
		.chanx_left_in(sb_1__1__330_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__349_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__364_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__364_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__1_ (
		.chanx_left_in(sb_1__1__331_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__350_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__365_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__365_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__2_ (
		.chanx_left_in(sb_1__1__332_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__351_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__366_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__366_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__3_ (
		.chanx_left_in(sb_1__1__333_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__352_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__367_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__367_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__6_ (
		.chanx_left_in(sb_1__1__334_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__353_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__368_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__368_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__7_ (
		.chanx_left_in(sb_1__1__335_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__354_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__369_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__369_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__8_ (
		.chanx_left_in(sb_1__1__336_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__355_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__370_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__370_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__9_ (
		.chanx_left_in(sb_1__1__337_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__356_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__371_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__371_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__10_ (
		.chanx_left_in(sb_1__1__338_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__357_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__372_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__372_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__11_ (
		.chanx_left_in(sb_1__1__339_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__358_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__373_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__373_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__12_ (
		.chanx_left_in(sb_1__1__340_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__359_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__374_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__374_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__13_ (
		.chanx_left_in(sb_1__1__341_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__360_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__375_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__375_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__14_ (
		.chanx_left_in(sb_1__1__342_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__361_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__376_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__376_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__15_ (
		.chanx_left_in(sb_1__1__343_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__362_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__377_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__377_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__16_ (
		.chanx_left_in(sb_1__1__344_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__363_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__378_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__378_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__17_ (
		.chanx_left_in(sb_1__1__345_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__364_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__379_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__379_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__18_ (
		.chanx_left_in(sb_1__1__346_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__365_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__380_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__380_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__19_ (
		.chanx_left_in(sb_1__1__347_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__366_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__381_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__381_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__20_ (
		.chanx_left_in(sb_1__1__348_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__367_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__382_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__382_chanx_right_out[0:228]));

	cbx_1__1_ cbx_21__21_ (
		.chanx_left_in(sb_1__1__349_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__1__368_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__383_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__383_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__1_ (
		.chanx_left_in(sb_1__1__350_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__0_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__384_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__384_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__2_ (
		.chanx_left_in(sb_1__1__351_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__1_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__385_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__385_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__3_ (
		.chanx_left_in(sb_1__1__352_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__2_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__386_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__386_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__6_ (
		.chanx_left_in(sb_1__1__353_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__3_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__387_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__387_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__7_ (
		.chanx_left_in(sb_1__1__354_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__4_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__388_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__388_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__8_ (
		.chanx_left_in(sb_1__1__355_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__5_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__389_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__389_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__9_ (
		.chanx_left_in(sb_1__1__356_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__6_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__390_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__390_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__10_ (
		.chanx_left_in(sb_1__1__357_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__7_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__391_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__391_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__11_ (
		.chanx_left_in(sb_1__1__358_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__8_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__392_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__392_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__12_ (
		.chanx_left_in(sb_1__1__359_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__9_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__393_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__393_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__13_ (
		.chanx_left_in(sb_1__1__360_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__10_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__394_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__394_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__14_ (
		.chanx_left_in(sb_1__1__361_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__11_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__395_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__395_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__15_ (
		.chanx_left_in(sb_1__1__362_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__12_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__396_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__396_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__16_ (
		.chanx_left_in(sb_1__1__363_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__13_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__397_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__397_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__17_ (
		.chanx_left_in(sb_1__1__364_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__14_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__398_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__398_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__18_ (
		.chanx_left_in(sb_1__1__365_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__15_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__399_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__399_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__19_ (
		.chanx_left_in(sb_1__1__366_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__16_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__400_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__400_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__20_ (
		.chanx_left_in(sb_1__1__367_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__17_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__401_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__401_chanx_right_out[0:228]));

	cbx_1__1_ cbx_22__21_ (
		.chanx_left_in(sb_1__1__368_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__1__18_chanx_left_out[0:228]),
		.chanx_left_out(cbx_1__1__402_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__1__402_chanx_right_out[0:228]));

	cbx_1__4_ cbx_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__4__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__0_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__0_ccff_tail),
		.chanx_left_out(cbx_1__4__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__0_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__0_ccff_tail));

	cbx_1__4_ cbx_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__1_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__1_ccff_tail),
		.chanx_left_out(cbx_1__4__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__1_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__1_ccff_tail));

	cbx_1__4_ cbx_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__2_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__2_ccff_tail),
		.chanx_left_out(cbx_1__4__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__2_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__2_ccff_tail));

	cbx_1__4_ cbx_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__3_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__3_ccff_tail),
		.chanx_left_out(cbx_1__4__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__3_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__3_ccff_tail));

	cbx_1__4_ cbx_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__4_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__4_ccff_tail),
		.chanx_left_out(cbx_1__4__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__4_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__4_ccff_tail));

	cbx_1__4_ cbx_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__5_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__5_ccff_tail),
		.chanx_left_out(cbx_1__4__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__5_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__5_ccff_tail));

	cbx_1__4_ cbx_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__6_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__6_ccff_tail),
		.chanx_left_out(cbx_1__4__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__6_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__6_ccff_tail));

	cbx_1__4_ cbx_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__7_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__7_ccff_tail),
		.chanx_left_out(cbx_1__4__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__7_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__7_ccff_tail));

	cbx_1__4_ cbx_9__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__8_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__8_ccff_tail),
		.chanx_left_out(cbx_1__4__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__8_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__8_ccff_tail));

	cbx_1__4_ cbx_10__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__9_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__9_ccff_tail),
		.chanx_left_out(cbx_1__4__9_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__9_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__9_ccff_tail));

	cbx_1__4_ cbx_11__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__10_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__10_ccff_tail),
		.chanx_left_out(cbx_1__4__10_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__10_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__10_ccff_tail));

	cbx_1__4_ cbx_12__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__11_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__11_ccff_tail),
		.chanx_left_out(cbx_1__4__11_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__11_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__11_ccff_tail));

	cbx_1__4_ cbx_13__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__12_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__12_ccff_tail),
		.chanx_left_out(cbx_1__4__12_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__12_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__12_ccff_tail));

	cbx_1__4_ cbx_14__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__13_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__13_ccff_tail),
		.chanx_left_out(cbx_1__4__13_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__13_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__13_ccff_tail));

	cbx_1__4_ cbx_15__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__14_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__14_ccff_tail),
		.chanx_left_out(cbx_1__4__14_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__14_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__14_ccff_tail));

	cbx_1__4_ cbx_16__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__15_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__15_ccff_tail),
		.chanx_left_out(cbx_1__4__15_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__15_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__15_ccff_tail));

	cbx_1__4_ cbx_17__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__15_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__16_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__16_ccff_tail),
		.chanx_left_out(cbx_1__4__16_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__16_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__16_ccff_tail));

	cbx_1__4_ cbx_18__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__16_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__17_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__17_ccff_tail),
		.chanx_left_out(cbx_1__4__17_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__17_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__17_ccff_tail));

	cbx_1__4_ cbx_19__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__17_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__18_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__18_ccff_tail),
		.chanx_left_out(cbx_1__4__18_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__18_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__18_ccff_tail));

	cbx_1__4_ cbx_20__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__18_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__19_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__19_ccff_tail),
		.chanx_left_out(cbx_1__4__19_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__19_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__19_ccff_tail));

	cbx_1__4_ cbx_21__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__19_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__4__20_chanx_left_out[0:228]),
		.ccff_head(sb_1__4__20_ccff_tail),
		.chanx_left_out(cbx_1__4__20_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__20_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__20_ccff_tail));

	cbx_1__4_ cbx_22__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__20_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__4__0_chanx_left_out[0:228]),
		.ccff_head(sb_22__4__0_ccff_tail),
		.chanx_left_out(cbx_1__4__21_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__4__21_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__4__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.ccff_tail(cbx_1__4__21_ccff_tail));

	cbx_1__5_ cbx_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__5__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__0_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__0_ccff_tail),
		.chanx_left_out(cbx_1__5__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__0_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__0_ccff_tail));

	cbx_1__5_ cbx_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__5__0_chanx_left_out[0:228]),
		.ccff_head(sb_2__5__0_ccff_tail),
		.chanx_left_out(cbx_1__5__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__1_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__1_ccff_tail));

	cbx_1__5_ cbx_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__5__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__1_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__1_ccff_tail),
		.chanx_left_out(cbx_1__5__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__2_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__2_ccff_tail));

	cbx_1__5_ cbx_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__5__1_chanx_left_out[0:228]),
		.ccff_head(sb_2__5__1_ccff_tail),
		.chanx_left_out(cbx_1__5__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__3_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__3_ccff_tail));

	cbx_1__5_ cbx_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__5__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__2_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__2_ccff_tail),
		.chanx_left_out(cbx_1__5__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__4_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__4_ccff_tail));

	cbx_1__5_ cbx_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_2__5__2_chanx_left_out[0:228]),
		.ccff_head(sb_2__5__2_ccff_tail),
		.chanx_left_out(cbx_1__5__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__5_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__5_ccff_tail));

	cbx_1__5_ cbx_10__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__5__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__3_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__3_ccff_tail),
		.chanx_left_out(cbx_1__5__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__6_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__6_ccff_tail));

	cbx_1__5_ cbx_11__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__4_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__4_ccff_tail),
		.chanx_left_out(cbx_1__5__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__7_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__7_ccff_tail));

	cbx_1__5_ cbx_12__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__5_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__5_ccff_tail),
		.chanx_left_out(cbx_1__5__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__8_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__8_ccff_tail));

	cbx_1__5_ cbx_13__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__6_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__6_ccff_tail),
		.chanx_left_out(cbx_1__5__9_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__9_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__9_ccff_tail));

	cbx_1__5_ cbx_14__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__7_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__7_ccff_tail),
		.chanx_left_out(cbx_1__5__10_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__10_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__10_ccff_tail));

	cbx_1__5_ cbx_15__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__8_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__8_ccff_tail),
		.chanx_left_out(cbx_1__5__11_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__11_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__11_ccff_tail));

	cbx_1__5_ cbx_16__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__9_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__9_ccff_tail),
		.chanx_left_out(cbx_1__5__12_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__12_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__12_ccff_tail));

	cbx_1__5_ cbx_17__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__10_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__10_ccff_tail),
		.chanx_left_out(cbx_1__5__13_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__13_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__13_ccff_tail));

	cbx_1__5_ cbx_18__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__11_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__11_ccff_tail),
		.chanx_left_out(cbx_1__5__14_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__14_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__14_ccff_tail));

	cbx_1__5_ cbx_19__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__12_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__12_ccff_tail),
		.chanx_left_out(cbx_1__5__15_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__15_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__15_ccff_tail));

	cbx_1__5_ cbx_20__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__13_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__13_ccff_tail),
		.chanx_left_out(cbx_1__5__16_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__16_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__16_ccff_tail));

	cbx_1__5_ cbx_21__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__5__14_chanx_left_out[0:228]),
		.ccff_head(sb_1__5__14_ccff_tail),
		.chanx_left_out(cbx_1__5__17_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__17_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__17_ccff_tail));

	cbx_1__5_ cbx_22__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__5__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__5__0_chanx_left_out[0:228]),
		.ccff_head(sb_22__5__0_ccff_tail),
		.chanx_left_out(cbx_1__5__18_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__5__18_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__5__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__5__18_ccff_tail));

	cbx_1__22_ cbx_1__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__22__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__0_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__0_ccff_tail),
		.chanx_left_out(cbx_1__22__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__0_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__0_ccff_tail));

	cbx_1__22_ cbx_2__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__1_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__1_ccff_tail),
		.chanx_left_out(cbx_1__22__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__1_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__1_ccff_tail));

	cbx_1__22_ cbx_3__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__2_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__2_ccff_tail),
		.chanx_left_out(cbx_1__22__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__2_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__2_ccff_tail));

	cbx_1__22_ cbx_4__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__3_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__3_ccff_tail),
		.chanx_left_out(cbx_1__22__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__3_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__3_ccff_tail));

	cbx_1__22_ cbx_5__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__4_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__4_ccff_tail),
		.chanx_left_out(cbx_1__22__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__4_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__4_ccff_tail));

	cbx_1__22_ cbx_6__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__5_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__5_ccff_tail),
		.chanx_left_out(cbx_1__22__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__5_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__5_ccff_tail));

	cbx_1__22_ cbx_7__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__6_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__6_ccff_tail),
		.chanx_left_out(cbx_1__22__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__6_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__6_ccff_tail));

	cbx_1__22_ cbx_8__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__7_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__7_ccff_tail),
		.chanx_left_out(cbx_1__22__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__7_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__7_ccff_tail));

	cbx_1__22_ cbx_9__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__8_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__8_ccff_tail),
		.chanx_left_out(cbx_1__22__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__8_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__8_ccff_tail));

	cbx_1__22_ cbx_10__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__9_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__9_ccff_tail),
		.chanx_left_out(cbx_1__22__9_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__9_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__9_ccff_tail));

	cbx_1__22_ cbx_11__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__9_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__10_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__10_ccff_tail),
		.chanx_left_out(cbx_1__22__10_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__10_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__10_ccff_tail));

	cbx_1__22_ cbx_12__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__10_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__11_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__11_ccff_tail),
		.chanx_left_out(cbx_1__22__11_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__11_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__11_ccff_tail));

	cbx_1__22_ cbx_13__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__11_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__12_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__12_ccff_tail),
		.chanx_left_out(cbx_1__22__12_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__12_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__12_ccff_tail));

	cbx_1__22_ cbx_14__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__12_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__13_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__13_ccff_tail),
		.chanx_left_out(cbx_1__22__13_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__13_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__13_ccff_tail));

	cbx_1__22_ cbx_15__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__13_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__14_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__14_ccff_tail),
		.chanx_left_out(cbx_1__22__14_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__14_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__14_ccff_tail));

	cbx_1__22_ cbx_16__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__14_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__15_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__15_ccff_tail),
		.chanx_left_out(cbx_1__22__15_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__15_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__15_ccff_tail));

	cbx_1__22_ cbx_17__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__15_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__16_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__16_ccff_tail),
		.chanx_left_out(cbx_1__22__16_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__16_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__16_ccff_tail));

	cbx_1__22_ cbx_18__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__16_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__17_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__17_ccff_tail),
		.chanx_left_out(cbx_1__22__17_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__17_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__17_ccff_tail));

	cbx_1__22_ cbx_19__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__17_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__18_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__18_ccff_tail),
		.chanx_left_out(cbx_1__22__18_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__18_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__18_ccff_tail));

	cbx_1__22_ cbx_20__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__18_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__19_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__19_ccff_tail),
		.chanx_left_out(cbx_1__22__19_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__19_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__19_ccff_tail));

	cbx_1__22_ cbx_21__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__19_chanx_right_out[0:228]),
		.chanx_right_in(sb_1__22__20_chanx_left_out[0:228]),
		.ccff_head(sb_1__22__20_ccff_tail),
		.chanx_left_out(cbx_1__22__20_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__20_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__20_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__20_ccff_tail));

	cbx_1__22_ cbx_22__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__22__20_chanx_right_out[0:228]),
		.chanx_right_in(sb_22__22__0_chanx_left_out[0:228]),
		.ccff_head(sb_22__22__0_ccff_tail),
		.chanx_left_out(cbx_1__22__21_chanx_left_out[0:228]),
		.chanx_right_out(cbx_1__22__21_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__22__21_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__22__21_ccff_tail));

	cbx_3__2_ cbx_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__0_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__0_ccff_tail),
		.chanx_left_out(cbx_3__2__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__0_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__0_ccff_tail));

	cbx_3__2_ cbx_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__1_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__1_ccff_tail),
		.chanx_left_out(cbx_3__2__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__1_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__1_ccff_tail));

	cbx_3__2_ cbx_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__2_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__2_ccff_tail),
		.chanx_left_out(cbx_3__2__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__2_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__2_ccff_tail));

	cbx_3__2_ cbx_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__3_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__3_ccff_tail),
		.chanx_left_out(cbx_3__2__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__3_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__3_ccff_tail));

	cbx_3__2_ cbx_9__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__4_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__4_ccff_tail),
		.chanx_left_out(cbx_3__2__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__4_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__4_ccff_tail));

	cbx_3__2_ cbx_9__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__2__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__2__5_chanx_left_out[0:228]),
		.ccff_head(sb_3__2__5_ccff_tail),
		.chanx_left_out(cbx_3__2__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__2__5_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.ccff_tail(cbx_3__2__5_ccff_tail));

	cbx_3__3_ cbx_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__0_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__0_ccff_tail),
		.chanx_left_out(cbx_3__3__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__0_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__0_ccff_tail));

	cbx_3__3_ cbx_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__1_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__1_ccff_tail),
		.chanx_left_out(cbx_3__3__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__1_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__1_ccff_tail));

	cbx_3__3_ cbx_3__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__2_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__2_ccff_tail),
		.chanx_left_out(cbx_3__3__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__2_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__2_ccff_tail));

	cbx_3__3_ cbx_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__3_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__3_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__3_ccff_tail),
		.chanx_left_out(cbx_3__3__3_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__3_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__3_ccff_tail));

	cbx_3__3_ cbx_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__4_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__4_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__4_ccff_tail),
		.chanx_left_out(cbx_3__3__4_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__4_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__4_ccff_tail));

	cbx_3__3_ cbx_6__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__5_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__5_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__5_ccff_tail),
		.chanx_left_out(cbx_3__3__5_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__5_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__5_ccff_tail));

	cbx_3__3_ cbx_9__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__6_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__6_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__6_ccff_tail),
		.chanx_left_out(cbx_3__3__6_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__6_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__6_ccff_tail));

	cbx_3__3_ cbx_9__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__7_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__7_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__7_ccff_tail),
		.chanx_left_out(cbx_3__3__7_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__7_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__7_ccff_tail));

	cbx_3__3_ cbx_9__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__3__8_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__3__8_chanx_left_out[0:228]),
		.ccff_head(sb_3__3__8_ccff_tail),
		.chanx_left_out(cbx_3__3__8_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__3__8_chanx_right_out[0:228]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_4_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_(cbx_3__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cbx_3__3__8_ccff_tail));

	cbx_3__5_ cbx_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__5__0_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__5__0_chanx_left_out[0:228]),
		.ccff_head(sb_3__5__0_ccff_tail),
		.chanx_left_out(cbx_3__5__0_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__5__0_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_3__5__0_ccff_tail));

	cbx_3__5_ cbx_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__5__1_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__5__1_chanx_left_out[0:228]),
		.ccff_head(sb_3__5__1_ccff_tail),
		.chanx_left_out(cbx_3__5__1_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__5__1_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_3__5__1_ccff_tail));

	cbx_3__5_ cbx_9__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_2__5__2_chanx_right_out[0:228]),
		.chanx_right_in(sb_3__5__2_chanx_left_out[0:228]),
		.ccff_head(sb_3__5__2_ccff_tail),
		.chanx_left_out(cbx_3__5__2_chanx_left_out[0:228]),
		.chanx_right_out(cbx_3__5__2_chanx_right_out[0:228]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_(cbx_3__5__2_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_3__5__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_3__5__2_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:228]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:228]),
		.chany_top_in(sb_0__4__0_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__5__0_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:228]),
		.ccff_head(sb_0__5__0_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__1_ cby_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__5_ccff_tail));

	cby_0__1_ cby_0__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__4_ccff_tail),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__6_ccff_tail));

	cby_0__1_ cby_0__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__5_ccff_tail),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__7_ccff_tail));

	cby_0__1_ cby_0__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__7_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__6_ccff_tail),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__8_ccff_tail));

	cby_0__1_ cby_0__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__7_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__8_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__7_ccff_tail),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__9_ccff_tail));

	cby_0__1_ cby_0__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__8_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__9_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__8_ccff_tail),
		.chany_bottom_out(cby_0__1__10_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__10_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__10_ccff_tail));

	cby_0__1_ cby_0__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__9_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__10_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__9_ccff_tail),
		.chany_bottom_out(cby_0__1__11_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__11_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__11_ccff_tail));

	cby_0__1_ cby_0__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__10_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__11_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__10_ccff_tail),
		.chany_bottom_out(cby_0__1__12_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__12_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__12_ccff_tail));

	cby_0__1_ cby_0__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__11_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__12_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__11_ccff_tail),
		.chany_bottom_out(cby_0__1__13_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__13_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__13_ccff_tail));

	cby_0__1_ cby_0__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__12_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__13_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__12_ccff_tail),
		.chany_bottom_out(cby_0__1__14_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__14_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__14_ccff_tail));

	cby_0__1_ cby_0__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__13_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__14_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__13_ccff_tail),
		.chany_bottom_out(cby_0__1__15_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__15_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__15_ccff_tail));

	cby_0__1_ cby_0__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__14_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__15_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__14_ccff_tail),
		.chany_bottom_out(cby_0__1__16_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__16_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__16_ccff_tail));

	cby_0__1_ cby_0__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__15_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__16_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__15_ccff_tail),
		.chany_bottom_out(cby_0__1__17_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__17_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__17_ccff_tail));

	cby_0__1_ cby_0__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__16_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__17_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__16_ccff_tail),
		.chany_bottom_out(cby_0__1__18_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__18_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__18_ccff_tail));

	cby_0__1_ cby_0__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__17_chany_top_out[0:228]),
		.chany_top_in(sb_0__1__18_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__17_ccff_tail),
		.chany_bottom_out(cby_0__1__19_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__19_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__19_ccff_tail));

	cby_0__1_ cby_0__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__18_chany_top_out[0:228]),
		.chany_top_in(sb_0__22__0_chany_bottom_out[0:228]),
		.ccff_head(sb_0__1__18_ccff_tail),
		.chany_bottom_out(cby_0__1__20_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__1__20_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__20_ccff_tail));

	cby_0__5_ cby_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__4__0_chany_top_out[0:228]),
		.chany_top_in(sb_0__5__0_chany_bottom_out[0:228]),
		.ccff_head(sb_0__4__0_ccff_tail),
		.chany_bottom_out(cby_0__5__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_0__5__0_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__5__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__5__0_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:228]));

	cby_1__1_ cby_1__2_ (
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:228]));

	cby_1__1_ cby_1__3_ (
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:228]));

	cby_1__1_ cby_1__4_ (
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__0_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:228]));

	cby_1__1_ cby_1__6_ (
		.chany_bottom_in(sb_1__5__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:228]));

	cby_1__1_ cby_1__7_ (
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:228]));

	cby_1__1_ cby_1__8_ (
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:228]));

	cby_1__1_ cby_1__9_ (
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:228]));

	cby_1__1_ cby_1__10_ (
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:228]));

	cby_1__1_ cby_1__11_ (
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:228]));

	cby_1__1_ cby_1__12_ (
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:228]));

	cby_1__1_ cby_1__13_ (
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:228]));

	cby_1__1_ cby_1__14_ (
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:228]));

	cby_1__1_ cby_1__15_ (
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:228]));

	cby_1__1_ cby_1__16_ (
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:228]));

	cby_1__1_ cby_1__17_ (
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:228]));

	cby_1__1_ cby_1__18_ (
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:228]));

	cby_1__1_ cby_1__19_ (
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:228]));

	cby_1__1_ cby_1__20_ (
		.chany_bottom_in(sb_1__1__16_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:228]));

	cby_1__1_ cby_1__21_ (
		.chany_bottom_in(sb_1__1__17_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:228]));

	cby_1__1_ cby_1__22_ (
		.chany_bottom_in(sb_1__1__18_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__0_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:228]));

	cby_1__1_ cby_2__1_ (
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:228]));

	cby_1__1_ cby_2__2_ (
		.chany_bottom_in(sb_1__1__19_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__0_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:228]));

	cby_1__1_ cby_2__4_ (
		.chany_bottom_in(sb_2__3__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__1_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:228]));

	cby_1__1_ cby_2__7_ (
		.chany_bottom_in(sb_2__3__1_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:228]));

	cby_1__1_ cby_2__8_ (
		.chany_bottom_in(sb_1__1__20_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__1_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:228]));

	cby_1__1_ cby_2__10_ (
		.chany_bottom_in(sb_2__3__2_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:228]));

	cby_1__1_ cby_2__11_ (
		.chany_bottom_in(sb_1__1__21_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:228]));

	cby_1__1_ cby_2__12_ (
		.chany_bottom_in(sb_1__1__22_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:228]));

	cby_1__1_ cby_2__13_ (
		.chany_bottom_in(sb_1__1__23_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:228]));

	cby_1__1_ cby_2__14_ (
		.chany_bottom_in(sb_1__1__24_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:228]));

	cby_1__1_ cby_2__15_ (
		.chany_bottom_in(sb_1__1__25_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:228]));

	cby_1__1_ cby_2__16_ (
		.chany_bottom_in(sb_1__1__26_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:228]));

	cby_1__1_ cby_2__17_ (
		.chany_bottom_in(sb_1__1__27_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:228]));

	cby_1__1_ cby_2__18_ (
		.chany_bottom_in(sb_1__1__28_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:228]));

	cby_1__1_ cby_2__19_ (
		.chany_bottom_in(sb_1__1__29_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:228]));

	cby_1__1_ cby_2__20_ (
		.chany_bottom_in(sb_1__1__30_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:228]));

	cby_1__1_ cby_2__21_ (
		.chany_bottom_in(sb_1__1__31_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:228]));

	cby_1__1_ cby_2__22_ (
		.chany_bottom_in(sb_1__1__32_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__1_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:228]));

	cby_1__1_ cby_3__1_ (
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:228]));

	cby_1__1_ cby_3__2_ (
		.chany_bottom_in(sb_1__1__33_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__0_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:228]));

	cby_1__1_ cby_3__4_ (
		.chany_bottom_in(sb_3__3__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__2_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:228]));

	cby_1__1_ cby_3__7_ (
		.chany_bottom_in(sb_3__3__1_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:228]));

	cby_1__1_ cby_3__8_ (
		.chany_bottom_in(sb_1__1__34_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__1_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:228]));

	cby_1__1_ cby_3__10_ (
		.chany_bottom_in(sb_3__3__2_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:228]));

	cby_1__1_ cby_3__11_ (
		.chany_bottom_in(sb_1__1__35_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:228]));

	cby_1__1_ cby_3__12_ (
		.chany_bottom_in(sb_1__1__36_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:228]));

	cby_1__1_ cby_3__13_ (
		.chany_bottom_in(sb_1__1__37_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:228]));

	cby_1__1_ cby_3__14_ (
		.chany_bottom_in(sb_1__1__38_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:228]));

	cby_1__1_ cby_3__15_ (
		.chany_bottom_in(sb_1__1__39_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:228]));

	cby_1__1_ cby_3__16_ (
		.chany_bottom_in(sb_1__1__40_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:228]));

	cby_1__1_ cby_3__17_ (
		.chany_bottom_in(sb_1__1__41_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:228]));

	cby_1__1_ cby_3__18_ (
		.chany_bottom_in(sb_1__1__42_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:228]));

	cby_1__1_ cby_3__19_ (
		.chany_bottom_in(sb_1__1__43_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:228]));

	cby_1__1_ cby_3__20_ (
		.chany_bottom_in(sb_1__1__44_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:228]));

	cby_1__1_ cby_3__21_ (
		.chany_bottom_in(sb_1__1__45_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:228]));

	cby_1__1_ cby_3__22_ (
		.chany_bottom_in(sb_1__1__46_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__2_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__56_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__56_chany_top_out[0:228]));

	cby_1__1_ cby_4__1_ (
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__57_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__57_chany_top_out[0:228]));

	cby_1__1_ cby_4__2_ (
		.chany_bottom_in(sb_1__1__47_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__58_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__58_chany_top_out[0:228]));

	cby_1__1_ cby_4__3_ (
		.chany_bottom_in(sb_1__1__48_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__49_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__59_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__59_chany_top_out[0:228]));

	cby_1__1_ cby_4__4_ (
		.chany_bottom_in(sb_1__1__49_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__3_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__60_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__60_chany_top_out[0:228]));

	cby_1__1_ cby_4__6_ (
		.chany_bottom_in(sb_1__5__1_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__50_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__61_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__61_chany_top_out[0:228]));

	cby_1__1_ cby_4__7_ (
		.chany_bottom_in(sb_1__1__50_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__51_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__62_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__62_chany_top_out[0:228]));

	cby_1__1_ cby_4__8_ (
		.chany_bottom_in(sb_1__1__51_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__52_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__63_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__63_chany_top_out[0:228]));

	cby_1__1_ cby_4__9_ (
		.chany_bottom_in(sb_1__1__52_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__53_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__64_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__64_chany_top_out[0:228]));

	cby_1__1_ cby_4__10_ (
		.chany_bottom_in(sb_1__1__53_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__54_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__65_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__65_chany_top_out[0:228]));

	cby_1__1_ cby_4__11_ (
		.chany_bottom_in(sb_1__1__54_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__55_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__66_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__66_chany_top_out[0:228]));

	cby_1__1_ cby_4__12_ (
		.chany_bottom_in(sb_1__1__55_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__56_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__67_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__67_chany_top_out[0:228]));

	cby_1__1_ cby_4__13_ (
		.chany_bottom_in(sb_1__1__56_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__57_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__68_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__68_chany_top_out[0:228]));

	cby_1__1_ cby_4__14_ (
		.chany_bottom_in(sb_1__1__57_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__58_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__69_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__69_chany_top_out[0:228]));

	cby_1__1_ cby_4__15_ (
		.chany_bottom_in(sb_1__1__58_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__59_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__70_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__70_chany_top_out[0:228]));

	cby_1__1_ cby_4__16_ (
		.chany_bottom_in(sb_1__1__59_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__60_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__71_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__71_chany_top_out[0:228]));

	cby_1__1_ cby_4__17_ (
		.chany_bottom_in(sb_1__1__60_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__61_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__72_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__72_chany_top_out[0:228]));

	cby_1__1_ cby_4__18_ (
		.chany_bottom_in(sb_1__1__61_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__62_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__73_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__73_chany_top_out[0:228]));

	cby_1__1_ cby_4__19_ (
		.chany_bottom_in(sb_1__1__62_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__63_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__74_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__74_chany_top_out[0:228]));

	cby_1__1_ cby_4__20_ (
		.chany_bottom_in(sb_1__1__63_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__64_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__75_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__75_chany_top_out[0:228]));

	cby_1__1_ cby_4__21_ (
		.chany_bottom_in(sb_1__1__64_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__65_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__76_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__76_chany_top_out[0:228]));

	cby_1__1_ cby_4__22_ (
		.chany_bottom_in(sb_1__1__65_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__3_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__77_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__77_chany_top_out[0:228]));

	cby_1__1_ cby_5__1_ (
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__66_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__78_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__78_chany_top_out[0:228]));

	cby_1__1_ cby_5__2_ (
		.chany_bottom_in(sb_1__1__66_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__2_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__79_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__79_chany_top_out[0:228]));

	cby_1__1_ cby_5__4_ (
		.chany_bottom_in(sb_2__3__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__4_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__80_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__80_chany_top_out[0:228]));

	cby_1__1_ cby_5__7_ (
		.chany_bottom_in(sb_2__3__4_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__67_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__81_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__81_chany_top_out[0:228]));

	cby_1__1_ cby_5__8_ (
		.chany_bottom_in(sb_1__1__67_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__3_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__82_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__82_chany_top_out[0:228]));

	cby_1__1_ cby_5__10_ (
		.chany_bottom_in(sb_2__3__5_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__68_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__83_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__83_chany_top_out[0:228]));

	cby_1__1_ cby_5__11_ (
		.chany_bottom_in(sb_1__1__68_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__69_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__84_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__84_chany_top_out[0:228]));

	cby_1__1_ cby_5__12_ (
		.chany_bottom_in(sb_1__1__69_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__70_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__85_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__85_chany_top_out[0:228]));

	cby_1__1_ cby_5__13_ (
		.chany_bottom_in(sb_1__1__70_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__71_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__86_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__86_chany_top_out[0:228]));

	cby_1__1_ cby_5__14_ (
		.chany_bottom_in(sb_1__1__71_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__72_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__87_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__87_chany_top_out[0:228]));

	cby_1__1_ cby_5__15_ (
		.chany_bottom_in(sb_1__1__72_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__73_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__88_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__88_chany_top_out[0:228]));

	cby_1__1_ cby_5__16_ (
		.chany_bottom_in(sb_1__1__73_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__74_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__89_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__89_chany_top_out[0:228]));

	cby_1__1_ cby_5__17_ (
		.chany_bottom_in(sb_1__1__74_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__75_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__90_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__90_chany_top_out[0:228]));

	cby_1__1_ cby_5__18_ (
		.chany_bottom_in(sb_1__1__75_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__76_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__91_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__91_chany_top_out[0:228]));

	cby_1__1_ cby_5__19_ (
		.chany_bottom_in(sb_1__1__76_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__77_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__92_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__92_chany_top_out[0:228]));

	cby_1__1_ cby_5__20_ (
		.chany_bottom_in(sb_1__1__77_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__78_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__93_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__93_chany_top_out[0:228]));

	cby_1__1_ cby_5__21_ (
		.chany_bottom_in(sb_1__1__78_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__79_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__94_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__94_chany_top_out[0:228]));

	cby_1__1_ cby_5__22_ (
		.chany_bottom_in(sb_1__1__79_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__4_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__95_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__95_chany_top_out[0:228]));

	cby_1__1_ cby_6__1_ (
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__80_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__96_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__96_chany_top_out[0:228]));

	cby_1__1_ cby_6__2_ (
		.chany_bottom_in(sb_1__1__80_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__2_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__97_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__97_chany_top_out[0:228]));

	cby_1__1_ cby_6__4_ (
		.chany_bottom_in(sb_3__3__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__5_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__98_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__98_chany_top_out[0:228]));

	cby_1__1_ cby_6__7_ (
		.chany_bottom_in(sb_3__3__4_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__81_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__99_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__99_chany_top_out[0:228]));

	cby_1__1_ cby_6__8_ (
		.chany_bottom_in(sb_1__1__81_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__3_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__100_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__100_chany_top_out[0:228]));

	cby_1__1_ cby_6__10_ (
		.chany_bottom_in(sb_3__3__5_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__82_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__101_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__101_chany_top_out[0:228]));

	cby_1__1_ cby_6__11_ (
		.chany_bottom_in(sb_1__1__82_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__83_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__102_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__102_chany_top_out[0:228]));

	cby_1__1_ cby_6__12_ (
		.chany_bottom_in(sb_1__1__83_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__84_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__103_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__103_chany_top_out[0:228]));

	cby_1__1_ cby_6__13_ (
		.chany_bottom_in(sb_1__1__84_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__85_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__104_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__104_chany_top_out[0:228]));

	cby_1__1_ cby_6__14_ (
		.chany_bottom_in(sb_1__1__85_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__86_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__105_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__105_chany_top_out[0:228]));

	cby_1__1_ cby_6__15_ (
		.chany_bottom_in(sb_1__1__86_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__87_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__106_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__106_chany_top_out[0:228]));

	cby_1__1_ cby_6__16_ (
		.chany_bottom_in(sb_1__1__87_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__88_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__107_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__107_chany_top_out[0:228]));

	cby_1__1_ cby_6__17_ (
		.chany_bottom_in(sb_1__1__88_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__89_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__108_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__108_chany_top_out[0:228]));

	cby_1__1_ cby_6__18_ (
		.chany_bottom_in(sb_1__1__89_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__90_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__109_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__109_chany_top_out[0:228]));

	cby_1__1_ cby_6__19_ (
		.chany_bottom_in(sb_1__1__90_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__91_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__110_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__110_chany_top_out[0:228]));

	cby_1__1_ cby_6__20_ (
		.chany_bottom_in(sb_1__1__91_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__92_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__111_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__111_chany_top_out[0:228]));

	cby_1__1_ cby_6__21_ (
		.chany_bottom_in(sb_1__1__92_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__93_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__112_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__112_chany_top_out[0:228]));

	cby_1__1_ cby_6__22_ (
		.chany_bottom_in(sb_1__1__93_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__5_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__113_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__113_chany_top_out[0:228]));

	cby_1__1_ cby_7__1_ (
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__94_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__114_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__114_chany_top_out[0:228]));

	cby_1__1_ cby_7__2_ (
		.chany_bottom_in(sb_1__1__94_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__95_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__115_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__115_chany_top_out[0:228]));

	cby_1__1_ cby_7__3_ (
		.chany_bottom_in(sb_1__1__95_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__96_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__116_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__116_chany_top_out[0:228]));

	cby_1__1_ cby_7__4_ (
		.chany_bottom_in(sb_1__1__96_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__6_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__117_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__117_chany_top_out[0:228]));

	cby_1__1_ cby_7__6_ (
		.chany_bottom_in(sb_1__5__2_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__97_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__118_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__118_chany_top_out[0:228]));

	cby_1__1_ cby_7__7_ (
		.chany_bottom_in(sb_1__1__97_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__98_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__119_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__119_chany_top_out[0:228]));

	cby_1__1_ cby_7__8_ (
		.chany_bottom_in(sb_1__1__98_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__99_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__120_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__120_chany_top_out[0:228]));

	cby_1__1_ cby_7__9_ (
		.chany_bottom_in(sb_1__1__99_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__100_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__121_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__121_chany_top_out[0:228]));

	cby_1__1_ cby_7__10_ (
		.chany_bottom_in(sb_1__1__100_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__101_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__122_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__122_chany_top_out[0:228]));

	cby_1__1_ cby_7__11_ (
		.chany_bottom_in(sb_1__1__101_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__102_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__123_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__123_chany_top_out[0:228]));

	cby_1__1_ cby_7__12_ (
		.chany_bottom_in(sb_1__1__102_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__103_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__124_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__124_chany_top_out[0:228]));

	cby_1__1_ cby_7__13_ (
		.chany_bottom_in(sb_1__1__103_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__104_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__125_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__125_chany_top_out[0:228]));

	cby_1__1_ cby_7__14_ (
		.chany_bottom_in(sb_1__1__104_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__105_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__126_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__126_chany_top_out[0:228]));

	cby_1__1_ cby_7__15_ (
		.chany_bottom_in(sb_1__1__105_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__106_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__127_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__127_chany_top_out[0:228]));

	cby_1__1_ cby_7__16_ (
		.chany_bottom_in(sb_1__1__106_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__107_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__128_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__128_chany_top_out[0:228]));

	cby_1__1_ cby_7__17_ (
		.chany_bottom_in(sb_1__1__107_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__108_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__129_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__129_chany_top_out[0:228]));

	cby_1__1_ cby_7__18_ (
		.chany_bottom_in(sb_1__1__108_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__109_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__130_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__130_chany_top_out[0:228]));

	cby_1__1_ cby_7__19_ (
		.chany_bottom_in(sb_1__1__109_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__110_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__131_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__131_chany_top_out[0:228]));

	cby_1__1_ cby_7__20_ (
		.chany_bottom_in(sb_1__1__110_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__111_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__132_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__132_chany_top_out[0:228]));

	cby_1__1_ cby_7__21_ (
		.chany_bottom_in(sb_1__1__111_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__112_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__133_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__133_chany_top_out[0:228]));

	cby_1__1_ cby_7__22_ (
		.chany_bottom_in(sb_1__1__112_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__6_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__134_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__134_chany_top_out[0:228]));

	cby_1__1_ cby_8__1_ (
		.chany_bottom_in(sb_1__0__7_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__113_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__135_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__135_chany_top_out[0:228]));

	cby_1__1_ cby_8__2_ (
		.chany_bottom_in(sb_1__1__113_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__4_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__136_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__136_chany_top_out[0:228]));

	cby_1__1_ cby_8__4_ (
		.chany_bottom_in(sb_2__3__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__7_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__137_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__137_chany_top_out[0:228]));

	cby_1__1_ cby_8__7_ (
		.chany_bottom_in(sb_2__3__7_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__114_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__138_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__138_chany_top_out[0:228]));

	cby_1__1_ cby_8__8_ (
		.chany_bottom_in(sb_1__1__114_chany_top_out[0:228]),
		.chany_top_in(sb_2__2__5_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__139_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__139_chany_top_out[0:228]));

	cby_1__1_ cby_8__10_ (
		.chany_bottom_in(sb_2__3__8_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__115_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__140_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__140_chany_top_out[0:228]));

	cby_1__1_ cby_8__11_ (
		.chany_bottom_in(sb_1__1__115_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__116_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__141_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__141_chany_top_out[0:228]));

	cby_1__1_ cby_8__12_ (
		.chany_bottom_in(sb_1__1__116_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__117_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__142_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__142_chany_top_out[0:228]));

	cby_1__1_ cby_8__13_ (
		.chany_bottom_in(sb_1__1__117_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__118_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__143_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__143_chany_top_out[0:228]));

	cby_1__1_ cby_8__14_ (
		.chany_bottom_in(sb_1__1__118_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__119_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__144_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__144_chany_top_out[0:228]));

	cby_1__1_ cby_8__15_ (
		.chany_bottom_in(sb_1__1__119_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__120_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__145_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__145_chany_top_out[0:228]));

	cby_1__1_ cby_8__16_ (
		.chany_bottom_in(sb_1__1__120_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__121_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__146_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__146_chany_top_out[0:228]));

	cby_1__1_ cby_8__17_ (
		.chany_bottom_in(sb_1__1__121_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__122_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__147_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__147_chany_top_out[0:228]));

	cby_1__1_ cby_8__18_ (
		.chany_bottom_in(sb_1__1__122_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__123_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__148_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__148_chany_top_out[0:228]));

	cby_1__1_ cby_8__19_ (
		.chany_bottom_in(sb_1__1__123_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__124_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__149_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__149_chany_top_out[0:228]));

	cby_1__1_ cby_8__20_ (
		.chany_bottom_in(sb_1__1__124_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__125_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__150_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__150_chany_top_out[0:228]));

	cby_1__1_ cby_8__21_ (
		.chany_bottom_in(sb_1__1__125_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__126_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__151_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__151_chany_top_out[0:228]));

	cby_1__1_ cby_8__22_ (
		.chany_bottom_in(sb_1__1__126_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__7_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__152_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__152_chany_top_out[0:228]));

	cby_1__1_ cby_9__1_ (
		.chany_bottom_in(sb_1__0__8_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__127_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__153_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__153_chany_top_out[0:228]));

	cby_1__1_ cby_9__2_ (
		.chany_bottom_in(sb_1__1__127_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__4_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__154_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__154_chany_top_out[0:228]));

	cby_1__1_ cby_9__4_ (
		.chany_bottom_in(sb_3__3__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__8_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__155_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__155_chany_top_out[0:228]));

	cby_1__1_ cby_9__7_ (
		.chany_bottom_in(sb_3__3__7_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__128_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__156_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__156_chany_top_out[0:228]));

	cby_1__1_ cby_9__8_ (
		.chany_bottom_in(sb_1__1__128_chany_top_out[0:228]),
		.chany_top_in(sb_3__2__5_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__157_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__157_chany_top_out[0:228]));

	cby_1__1_ cby_9__10_ (
		.chany_bottom_in(sb_3__3__8_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__129_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__158_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__158_chany_top_out[0:228]));

	cby_1__1_ cby_9__11_ (
		.chany_bottom_in(sb_1__1__129_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__130_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__159_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__159_chany_top_out[0:228]));

	cby_1__1_ cby_9__12_ (
		.chany_bottom_in(sb_1__1__130_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__131_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__160_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__160_chany_top_out[0:228]));

	cby_1__1_ cby_9__13_ (
		.chany_bottom_in(sb_1__1__131_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__132_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__161_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__161_chany_top_out[0:228]));

	cby_1__1_ cby_9__14_ (
		.chany_bottom_in(sb_1__1__132_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__133_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__162_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__162_chany_top_out[0:228]));

	cby_1__1_ cby_9__15_ (
		.chany_bottom_in(sb_1__1__133_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__134_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__163_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__163_chany_top_out[0:228]));

	cby_1__1_ cby_9__16_ (
		.chany_bottom_in(sb_1__1__134_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__135_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__164_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__164_chany_top_out[0:228]));

	cby_1__1_ cby_9__17_ (
		.chany_bottom_in(sb_1__1__135_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__136_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__165_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__165_chany_top_out[0:228]));

	cby_1__1_ cby_9__18_ (
		.chany_bottom_in(sb_1__1__136_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__137_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__166_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__166_chany_top_out[0:228]));

	cby_1__1_ cby_9__19_ (
		.chany_bottom_in(sb_1__1__137_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__138_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__167_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__167_chany_top_out[0:228]));

	cby_1__1_ cby_9__20_ (
		.chany_bottom_in(sb_1__1__138_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__139_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__168_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__168_chany_top_out[0:228]));

	cby_1__1_ cby_9__21_ (
		.chany_bottom_in(sb_1__1__139_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__140_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__169_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__169_chany_top_out[0:228]));

	cby_1__1_ cby_9__22_ (
		.chany_bottom_in(sb_1__1__140_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__8_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__170_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__170_chany_top_out[0:228]));

	cby_1__1_ cby_10__1_ (
		.chany_bottom_in(sb_1__0__9_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__141_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__171_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__171_chany_top_out[0:228]));

	cby_1__1_ cby_10__2_ (
		.chany_bottom_in(sb_1__1__141_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__142_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__172_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__172_chany_top_out[0:228]));

	cby_1__1_ cby_10__3_ (
		.chany_bottom_in(sb_1__1__142_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__143_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__173_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__173_chany_top_out[0:228]));

	cby_1__1_ cby_10__4_ (
		.chany_bottom_in(sb_1__1__143_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__9_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__174_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__174_chany_top_out[0:228]));

	cby_1__1_ cby_10__6_ (
		.chany_bottom_in(sb_1__5__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__144_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__175_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__175_chany_top_out[0:228]));

	cby_1__1_ cby_10__7_ (
		.chany_bottom_in(sb_1__1__144_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__145_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__176_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__176_chany_top_out[0:228]));

	cby_1__1_ cby_10__8_ (
		.chany_bottom_in(sb_1__1__145_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__146_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__177_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__177_chany_top_out[0:228]));

	cby_1__1_ cby_10__9_ (
		.chany_bottom_in(sb_1__1__146_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__147_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__178_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__178_chany_top_out[0:228]));

	cby_1__1_ cby_10__10_ (
		.chany_bottom_in(sb_1__1__147_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__148_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__179_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__179_chany_top_out[0:228]));

	cby_1__1_ cby_10__11_ (
		.chany_bottom_in(sb_1__1__148_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__149_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__180_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__180_chany_top_out[0:228]));

	cby_1__1_ cby_10__12_ (
		.chany_bottom_in(sb_1__1__149_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__150_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__181_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__181_chany_top_out[0:228]));

	cby_1__1_ cby_10__13_ (
		.chany_bottom_in(sb_1__1__150_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__151_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__182_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__182_chany_top_out[0:228]));

	cby_1__1_ cby_10__14_ (
		.chany_bottom_in(sb_1__1__151_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__152_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__183_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__183_chany_top_out[0:228]));

	cby_1__1_ cby_10__15_ (
		.chany_bottom_in(sb_1__1__152_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__153_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__184_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__184_chany_top_out[0:228]));

	cby_1__1_ cby_10__16_ (
		.chany_bottom_in(sb_1__1__153_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__154_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__185_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__185_chany_top_out[0:228]));

	cby_1__1_ cby_10__17_ (
		.chany_bottom_in(sb_1__1__154_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__155_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__186_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__186_chany_top_out[0:228]));

	cby_1__1_ cby_10__18_ (
		.chany_bottom_in(sb_1__1__155_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__156_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__187_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__187_chany_top_out[0:228]));

	cby_1__1_ cby_10__19_ (
		.chany_bottom_in(sb_1__1__156_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__157_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__188_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__188_chany_top_out[0:228]));

	cby_1__1_ cby_10__20_ (
		.chany_bottom_in(sb_1__1__157_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__158_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__189_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__189_chany_top_out[0:228]));

	cby_1__1_ cby_10__21_ (
		.chany_bottom_in(sb_1__1__158_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__159_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__190_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__190_chany_top_out[0:228]));

	cby_1__1_ cby_10__22_ (
		.chany_bottom_in(sb_1__1__159_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__9_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__191_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__191_chany_top_out[0:228]));

	cby_1__1_ cby_11__1_ (
		.chany_bottom_in(sb_1__0__10_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__160_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__192_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__192_chany_top_out[0:228]));

	cby_1__1_ cby_11__2_ (
		.chany_bottom_in(sb_1__1__160_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__161_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__193_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__193_chany_top_out[0:228]));

	cby_1__1_ cby_11__3_ (
		.chany_bottom_in(sb_1__1__161_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__162_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__194_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__194_chany_top_out[0:228]));

	cby_1__1_ cby_11__4_ (
		.chany_bottom_in(sb_1__1__162_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__10_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__195_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__195_chany_top_out[0:228]));

	cby_1__1_ cby_11__6_ (
		.chany_bottom_in(sb_1__5__4_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__163_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__196_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__196_chany_top_out[0:228]));

	cby_1__1_ cby_11__7_ (
		.chany_bottom_in(sb_1__1__163_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__164_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__197_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__197_chany_top_out[0:228]));

	cby_1__1_ cby_11__8_ (
		.chany_bottom_in(sb_1__1__164_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__165_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__198_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__198_chany_top_out[0:228]));

	cby_1__1_ cby_11__9_ (
		.chany_bottom_in(sb_1__1__165_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__166_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__199_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__199_chany_top_out[0:228]));

	cby_1__1_ cby_11__10_ (
		.chany_bottom_in(sb_1__1__166_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__167_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__200_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__200_chany_top_out[0:228]));

	cby_1__1_ cby_11__11_ (
		.chany_bottom_in(sb_1__1__167_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__168_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__201_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__201_chany_top_out[0:228]));

	cby_1__1_ cby_11__12_ (
		.chany_bottom_in(sb_1__1__168_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__169_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__202_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__202_chany_top_out[0:228]));

	cby_1__1_ cby_11__13_ (
		.chany_bottom_in(sb_1__1__169_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__170_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__203_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__203_chany_top_out[0:228]));

	cby_1__1_ cby_11__14_ (
		.chany_bottom_in(sb_1__1__170_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__171_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__204_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__204_chany_top_out[0:228]));

	cby_1__1_ cby_11__15_ (
		.chany_bottom_in(sb_1__1__171_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__172_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__205_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__205_chany_top_out[0:228]));

	cby_1__1_ cby_11__16_ (
		.chany_bottom_in(sb_1__1__172_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__173_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__206_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__206_chany_top_out[0:228]));

	cby_1__1_ cby_11__17_ (
		.chany_bottom_in(sb_1__1__173_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__174_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__207_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__207_chany_top_out[0:228]));

	cby_1__1_ cby_11__18_ (
		.chany_bottom_in(sb_1__1__174_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__175_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__208_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__208_chany_top_out[0:228]));

	cby_1__1_ cby_11__19_ (
		.chany_bottom_in(sb_1__1__175_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__176_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__209_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__209_chany_top_out[0:228]));

	cby_1__1_ cby_11__20_ (
		.chany_bottom_in(sb_1__1__176_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__177_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__210_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__210_chany_top_out[0:228]));

	cby_1__1_ cby_11__21_ (
		.chany_bottom_in(sb_1__1__177_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__178_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__211_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__211_chany_top_out[0:228]));

	cby_1__1_ cby_11__22_ (
		.chany_bottom_in(sb_1__1__178_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__10_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__212_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__212_chany_top_out[0:228]));

	cby_1__1_ cby_12__1_ (
		.chany_bottom_in(sb_1__0__11_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__179_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__213_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__213_chany_top_out[0:228]));

	cby_1__1_ cby_12__2_ (
		.chany_bottom_in(sb_1__1__179_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__180_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__214_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__214_chany_top_out[0:228]));

	cby_1__1_ cby_12__3_ (
		.chany_bottom_in(sb_1__1__180_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__181_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__215_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__215_chany_top_out[0:228]));

	cby_1__1_ cby_12__4_ (
		.chany_bottom_in(sb_1__1__181_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__11_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__216_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__216_chany_top_out[0:228]));

	cby_1__1_ cby_12__6_ (
		.chany_bottom_in(sb_1__5__5_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__182_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__217_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__217_chany_top_out[0:228]));

	cby_1__1_ cby_12__7_ (
		.chany_bottom_in(sb_1__1__182_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__183_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__218_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__218_chany_top_out[0:228]));

	cby_1__1_ cby_12__8_ (
		.chany_bottom_in(sb_1__1__183_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__184_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__219_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__219_chany_top_out[0:228]));

	cby_1__1_ cby_12__9_ (
		.chany_bottom_in(sb_1__1__184_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__185_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__220_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__220_chany_top_out[0:228]));

	cby_1__1_ cby_12__10_ (
		.chany_bottom_in(sb_1__1__185_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__186_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__221_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__221_chany_top_out[0:228]));

	cby_1__1_ cby_12__11_ (
		.chany_bottom_in(sb_1__1__186_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__187_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__222_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__222_chany_top_out[0:228]));

	cby_1__1_ cby_12__12_ (
		.chany_bottom_in(sb_1__1__187_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__188_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__223_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__223_chany_top_out[0:228]));

	cby_1__1_ cby_12__13_ (
		.chany_bottom_in(sb_1__1__188_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__189_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__224_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__224_chany_top_out[0:228]));

	cby_1__1_ cby_12__14_ (
		.chany_bottom_in(sb_1__1__189_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__190_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__225_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__225_chany_top_out[0:228]));

	cby_1__1_ cby_12__15_ (
		.chany_bottom_in(sb_1__1__190_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__191_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__226_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__226_chany_top_out[0:228]));

	cby_1__1_ cby_12__16_ (
		.chany_bottom_in(sb_1__1__191_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__192_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__227_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__227_chany_top_out[0:228]));

	cby_1__1_ cby_12__17_ (
		.chany_bottom_in(sb_1__1__192_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__193_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__228_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__228_chany_top_out[0:228]));

	cby_1__1_ cby_12__18_ (
		.chany_bottom_in(sb_1__1__193_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__194_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__229_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__229_chany_top_out[0:228]));

	cby_1__1_ cby_12__19_ (
		.chany_bottom_in(sb_1__1__194_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__195_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__230_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__230_chany_top_out[0:228]));

	cby_1__1_ cby_12__20_ (
		.chany_bottom_in(sb_1__1__195_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__196_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__231_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__231_chany_top_out[0:228]));

	cby_1__1_ cby_12__21_ (
		.chany_bottom_in(sb_1__1__196_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__197_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__232_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__232_chany_top_out[0:228]));

	cby_1__1_ cby_12__22_ (
		.chany_bottom_in(sb_1__1__197_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__11_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__233_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__233_chany_top_out[0:228]));

	cby_1__1_ cby_13__1_ (
		.chany_bottom_in(sb_1__0__12_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__198_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__234_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__234_chany_top_out[0:228]));

	cby_1__1_ cby_13__2_ (
		.chany_bottom_in(sb_1__1__198_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__199_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__235_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__235_chany_top_out[0:228]));

	cby_1__1_ cby_13__3_ (
		.chany_bottom_in(sb_1__1__199_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__200_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__236_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__236_chany_top_out[0:228]));

	cby_1__1_ cby_13__4_ (
		.chany_bottom_in(sb_1__1__200_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__12_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__237_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__237_chany_top_out[0:228]));

	cby_1__1_ cby_13__6_ (
		.chany_bottom_in(sb_1__5__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__201_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__238_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__238_chany_top_out[0:228]));

	cby_1__1_ cby_13__7_ (
		.chany_bottom_in(sb_1__1__201_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__202_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__239_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__239_chany_top_out[0:228]));

	cby_1__1_ cby_13__8_ (
		.chany_bottom_in(sb_1__1__202_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__203_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__240_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__240_chany_top_out[0:228]));

	cby_1__1_ cby_13__9_ (
		.chany_bottom_in(sb_1__1__203_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__204_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__241_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__241_chany_top_out[0:228]));

	cby_1__1_ cby_13__10_ (
		.chany_bottom_in(sb_1__1__204_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__205_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__242_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__242_chany_top_out[0:228]));

	cby_1__1_ cby_13__11_ (
		.chany_bottom_in(sb_1__1__205_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__206_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__243_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__243_chany_top_out[0:228]));

	cby_1__1_ cby_13__12_ (
		.chany_bottom_in(sb_1__1__206_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__207_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__244_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__244_chany_top_out[0:228]));

	cby_1__1_ cby_13__13_ (
		.chany_bottom_in(sb_1__1__207_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__208_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__245_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__245_chany_top_out[0:228]));

	cby_1__1_ cby_13__14_ (
		.chany_bottom_in(sb_1__1__208_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__209_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__246_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__246_chany_top_out[0:228]));

	cby_1__1_ cby_13__15_ (
		.chany_bottom_in(sb_1__1__209_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__210_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__247_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__247_chany_top_out[0:228]));

	cby_1__1_ cby_13__16_ (
		.chany_bottom_in(sb_1__1__210_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__211_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__248_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__248_chany_top_out[0:228]));

	cby_1__1_ cby_13__17_ (
		.chany_bottom_in(sb_1__1__211_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__212_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__249_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__249_chany_top_out[0:228]));

	cby_1__1_ cby_13__18_ (
		.chany_bottom_in(sb_1__1__212_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__213_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__250_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__250_chany_top_out[0:228]));

	cby_1__1_ cby_13__19_ (
		.chany_bottom_in(sb_1__1__213_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__214_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__251_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__251_chany_top_out[0:228]));

	cby_1__1_ cby_13__20_ (
		.chany_bottom_in(sb_1__1__214_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__215_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__252_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__252_chany_top_out[0:228]));

	cby_1__1_ cby_13__21_ (
		.chany_bottom_in(sb_1__1__215_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__216_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__253_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__253_chany_top_out[0:228]));

	cby_1__1_ cby_13__22_ (
		.chany_bottom_in(sb_1__1__216_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__12_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__254_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__254_chany_top_out[0:228]));

	cby_1__1_ cby_14__1_ (
		.chany_bottom_in(sb_1__0__13_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__217_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__255_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__255_chany_top_out[0:228]));

	cby_1__1_ cby_14__2_ (
		.chany_bottom_in(sb_1__1__217_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__218_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__256_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__256_chany_top_out[0:228]));

	cby_1__1_ cby_14__3_ (
		.chany_bottom_in(sb_1__1__218_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__219_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__257_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__257_chany_top_out[0:228]));

	cby_1__1_ cby_14__4_ (
		.chany_bottom_in(sb_1__1__219_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__13_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__258_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__258_chany_top_out[0:228]));

	cby_1__1_ cby_14__6_ (
		.chany_bottom_in(sb_1__5__7_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__220_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__259_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__259_chany_top_out[0:228]));

	cby_1__1_ cby_14__7_ (
		.chany_bottom_in(sb_1__1__220_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__221_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__260_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__260_chany_top_out[0:228]));

	cby_1__1_ cby_14__8_ (
		.chany_bottom_in(sb_1__1__221_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__222_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__261_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__261_chany_top_out[0:228]));

	cby_1__1_ cby_14__9_ (
		.chany_bottom_in(sb_1__1__222_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__223_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__262_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__262_chany_top_out[0:228]));

	cby_1__1_ cby_14__10_ (
		.chany_bottom_in(sb_1__1__223_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__224_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__263_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__263_chany_top_out[0:228]));

	cby_1__1_ cby_14__11_ (
		.chany_bottom_in(sb_1__1__224_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__225_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__264_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__264_chany_top_out[0:228]));

	cby_1__1_ cby_14__12_ (
		.chany_bottom_in(sb_1__1__225_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__226_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__265_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__265_chany_top_out[0:228]));

	cby_1__1_ cby_14__13_ (
		.chany_bottom_in(sb_1__1__226_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__227_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__266_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__266_chany_top_out[0:228]));

	cby_1__1_ cby_14__14_ (
		.chany_bottom_in(sb_1__1__227_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__228_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__267_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__267_chany_top_out[0:228]));

	cby_1__1_ cby_14__15_ (
		.chany_bottom_in(sb_1__1__228_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__229_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__268_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__268_chany_top_out[0:228]));

	cby_1__1_ cby_14__16_ (
		.chany_bottom_in(sb_1__1__229_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__230_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__269_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__269_chany_top_out[0:228]));

	cby_1__1_ cby_14__17_ (
		.chany_bottom_in(sb_1__1__230_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__231_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__270_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__270_chany_top_out[0:228]));

	cby_1__1_ cby_14__18_ (
		.chany_bottom_in(sb_1__1__231_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__232_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__271_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__271_chany_top_out[0:228]));

	cby_1__1_ cby_14__19_ (
		.chany_bottom_in(sb_1__1__232_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__233_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__272_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__272_chany_top_out[0:228]));

	cby_1__1_ cby_14__20_ (
		.chany_bottom_in(sb_1__1__233_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__234_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__273_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__273_chany_top_out[0:228]));

	cby_1__1_ cby_14__21_ (
		.chany_bottom_in(sb_1__1__234_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__235_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__274_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__274_chany_top_out[0:228]));

	cby_1__1_ cby_14__22_ (
		.chany_bottom_in(sb_1__1__235_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__13_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__275_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__275_chany_top_out[0:228]));

	cby_1__1_ cby_15__1_ (
		.chany_bottom_in(sb_1__0__14_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__236_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__276_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__276_chany_top_out[0:228]));

	cby_1__1_ cby_15__2_ (
		.chany_bottom_in(sb_1__1__236_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__237_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__277_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__277_chany_top_out[0:228]));

	cby_1__1_ cby_15__3_ (
		.chany_bottom_in(sb_1__1__237_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__238_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__278_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__278_chany_top_out[0:228]));

	cby_1__1_ cby_15__4_ (
		.chany_bottom_in(sb_1__1__238_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__14_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__279_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__279_chany_top_out[0:228]));

	cby_1__1_ cby_15__6_ (
		.chany_bottom_in(sb_1__5__8_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__239_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__280_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__280_chany_top_out[0:228]));

	cby_1__1_ cby_15__7_ (
		.chany_bottom_in(sb_1__1__239_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__240_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__281_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__281_chany_top_out[0:228]));

	cby_1__1_ cby_15__8_ (
		.chany_bottom_in(sb_1__1__240_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__241_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__282_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__282_chany_top_out[0:228]));

	cby_1__1_ cby_15__9_ (
		.chany_bottom_in(sb_1__1__241_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__242_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__283_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__283_chany_top_out[0:228]));

	cby_1__1_ cby_15__10_ (
		.chany_bottom_in(sb_1__1__242_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__243_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__284_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__284_chany_top_out[0:228]));

	cby_1__1_ cby_15__11_ (
		.chany_bottom_in(sb_1__1__243_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__244_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__285_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__285_chany_top_out[0:228]));

	cby_1__1_ cby_15__12_ (
		.chany_bottom_in(sb_1__1__244_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__245_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__286_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__286_chany_top_out[0:228]));

	cby_1__1_ cby_15__13_ (
		.chany_bottom_in(sb_1__1__245_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__246_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__287_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__287_chany_top_out[0:228]));

	cby_1__1_ cby_15__14_ (
		.chany_bottom_in(sb_1__1__246_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__247_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__288_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__288_chany_top_out[0:228]));

	cby_1__1_ cby_15__15_ (
		.chany_bottom_in(sb_1__1__247_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__248_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__289_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__289_chany_top_out[0:228]));

	cby_1__1_ cby_15__16_ (
		.chany_bottom_in(sb_1__1__248_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__249_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__290_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__290_chany_top_out[0:228]));

	cby_1__1_ cby_15__17_ (
		.chany_bottom_in(sb_1__1__249_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__250_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__291_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__291_chany_top_out[0:228]));

	cby_1__1_ cby_15__18_ (
		.chany_bottom_in(sb_1__1__250_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__251_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__292_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__292_chany_top_out[0:228]));

	cby_1__1_ cby_15__19_ (
		.chany_bottom_in(sb_1__1__251_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__252_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__293_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__293_chany_top_out[0:228]));

	cby_1__1_ cby_15__20_ (
		.chany_bottom_in(sb_1__1__252_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__253_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__294_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__294_chany_top_out[0:228]));

	cby_1__1_ cby_15__21_ (
		.chany_bottom_in(sb_1__1__253_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__254_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__295_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__295_chany_top_out[0:228]));

	cby_1__1_ cby_15__22_ (
		.chany_bottom_in(sb_1__1__254_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__14_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__296_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__296_chany_top_out[0:228]));

	cby_1__1_ cby_16__1_ (
		.chany_bottom_in(sb_1__0__15_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__255_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__297_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__297_chany_top_out[0:228]));

	cby_1__1_ cby_16__2_ (
		.chany_bottom_in(sb_1__1__255_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__256_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__298_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__298_chany_top_out[0:228]));

	cby_1__1_ cby_16__3_ (
		.chany_bottom_in(sb_1__1__256_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__257_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__299_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__299_chany_top_out[0:228]));

	cby_1__1_ cby_16__4_ (
		.chany_bottom_in(sb_1__1__257_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__15_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__300_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__300_chany_top_out[0:228]));

	cby_1__1_ cby_16__6_ (
		.chany_bottom_in(sb_1__5__9_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__258_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__301_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__301_chany_top_out[0:228]));

	cby_1__1_ cby_16__7_ (
		.chany_bottom_in(sb_1__1__258_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__259_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__302_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__302_chany_top_out[0:228]));

	cby_1__1_ cby_16__8_ (
		.chany_bottom_in(sb_1__1__259_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__260_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__303_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__303_chany_top_out[0:228]));

	cby_1__1_ cby_16__9_ (
		.chany_bottom_in(sb_1__1__260_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__261_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__304_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__304_chany_top_out[0:228]));

	cby_1__1_ cby_16__10_ (
		.chany_bottom_in(sb_1__1__261_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__262_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__305_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__305_chany_top_out[0:228]));

	cby_1__1_ cby_16__11_ (
		.chany_bottom_in(sb_1__1__262_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__263_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__306_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__306_chany_top_out[0:228]));

	cby_1__1_ cby_16__12_ (
		.chany_bottom_in(sb_1__1__263_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__264_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__307_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__307_chany_top_out[0:228]));

	cby_1__1_ cby_16__13_ (
		.chany_bottom_in(sb_1__1__264_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__265_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__308_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__308_chany_top_out[0:228]));

	cby_1__1_ cby_16__14_ (
		.chany_bottom_in(sb_1__1__265_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__266_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__309_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__309_chany_top_out[0:228]));

	cby_1__1_ cby_16__15_ (
		.chany_bottom_in(sb_1__1__266_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__267_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__310_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__310_chany_top_out[0:228]));

	cby_1__1_ cby_16__16_ (
		.chany_bottom_in(sb_1__1__267_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__268_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__311_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__311_chany_top_out[0:228]));

	cby_1__1_ cby_16__17_ (
		.chany_bottom_in(sb_1__1__268_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__269_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__312_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__312_chany_top_out[0:228]));

	cby_1__1_ cby_16__18_ (
		.chany_bottom_in(sb_1__1__269_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__270_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__313_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__313_chany_top_out[0:228]));

	cby_1__1_ cby_16__19_ (
		.chany_bottom_in(sb_1__1__270_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__271_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__314_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__314_chany_top_out[0:228]));

	cby_1__1_ cby_16__20_ (
		.chany_bottom_in(sb_1__1__271_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__272_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__315_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__315_chany_top_out[0:228]));

	cby_1__1_ cby_16__21_ (
		.chany_bottom_in(sb_1__1__272_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__273_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__316_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__316_chany_top_out[0:228]));

	cby_1__1_ cby_16__22_ (
		.chany_bottom_in(sb_1__1__273_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__15_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__317_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__317_chany_top_out[0:228]));

	cby_1__1_ cby_17__1_ (
		.chany_bottom_in(sb_1__0__16_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__274_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__318_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__318_chany_top_out[0:228]));

	cby_1__1_ cby_17__2_ (
		.chany_bottom_in(sb_1__1__274_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__275_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__319_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__319_chany_top_out[0:228]));

	cby_1__1_ cby_17__3_ (
		.chany_bottom_in(sb_1__1__275_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__276_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__320_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__320_chany_top_out[0:228]));

	cby_1__1_ cby_17__4_ (
		.chany_bottom_in(sb_1__1__276_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__16_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__321_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__321_chany_top_out[0:228]));

	cby_1__1_ cby_17__6_ (
		.chany_bottom_in(sb_1__5__10_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__277_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__322_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__322_chany_top_out[0:228]));

	cby_1__1_ cby_17__7_ (
		.chany_bottom_in(sb_1__1__277_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__278_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__323_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__323_chany_top_out[0:228]));

	cby_1__1_ cby_17__8_ (
		.chany_bottom_in(sb_1__1__278_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__279_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__324_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__324_chany_top_out[0:228]));

	cby_1__1_ cby_17__9_ (
		.chany_bottom_in(sb_1__1__279_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__280_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__325_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__325_chany_top_out[0:228]));

	cby_1__1_ cby_17__10_ (
		.chany_bottom_in(sb_1__1__280_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__281_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__326_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__326_chany_top_out[0:228]));

	cby_1__1_ cby_17__11_ (
		.chany_bottom_in(sb_1__1__281_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__282_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__327_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__327_chany_top_out[0:228]));

	cby_1__1_ cby_17__12_ (
		.chany_bottom_in(sb_1__1__282_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__283_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__328_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__328_chany_top_out[0:228]));

	cby_1__1_ cby_17__13_ (
		.chany_bottom_in(sb_1__1__283_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__284_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__329_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__329_chany_top_out[0:228]));

	cby_1__1_ cby_17__14_ (
		.chany_bottom_in(sb_1__1__284_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__285_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__330_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__330_chany_top_out[0:228]));

	cby_1__1_ cby_17__15_ (
		.chany_bottom_in(sb_1__1__285_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__286_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__331_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__331_chany_top_out[0:228]));

	cby_1__1_ cby_17__16_ (
		.chany_bottom_in(sb_1__1__286_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__287_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__332_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__332_chany_top_out[0:228]));

	cby_1__1_ cby_17__17_ (
		.chany_bottom_in(sb_1__1__287_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__288_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__333_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__333_chany_top_out[0:228]));

	cby_1__1_ cby_17__18_ (
		.chany_bottom_in(sb_1__1__288_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__289_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__334_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__334_chany_top_out[0:228]));

	cby_1__1_ cby_17__19_ (
		.chany_bottom_in(sb_1__1__289_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__290_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__335_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__335_chany_top_out[0:228]));

	cby_1__1_ cby_17__20_ (
		.chany_bottom_in(sb_1__1__290_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__291_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__336_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__336_chany_top_out[0:228]));

	cby_1__1_ cby_17__21_ (
		.chany_bottom_in(sb_1__1__291_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__292_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__337_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__337_chany_top_out[0:228]));

	cby_1__1_ cby_17__22_ (
		.chany_bottom_in(sb_1__1__292_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__16_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__338_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__338_chany_top_out[0:228]));

	cby_1__1_ cby_18__1_ (
		.chany_bottom_in(sb_1__0__17_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__293_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__339_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__339_chany_top_out[0:228]));

	cby_1__1_ cby_18__2_ (
		.chany_bottom_in(sb_1__1__293_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__294_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__340_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__340_chany_top_out[0:228]));

	cby_1__1_ cby_18__3_ (
		.chany_bottom_in(sb_1__1__294_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__295_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__341_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__341_chany_top_out[0:228]));

	cby_1__1_ cby_18__4_ (
		.chany_bottom_in(sb_1__1__295_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__17_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__342_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__342_chany_top_out[0:228]));

	cby_1__1_ cby_18__6_ (
		.chany_bottom_in(sb_1__5__11_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__296_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__343_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__343_chany_top_out[0:228]));

	cby_1__1_ cby_18__7_ (
		.chany_bottom_in(sb_1__1__296_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__297_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__344_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__344_chany_top_out[0:228]));

	cby_1__1_ cby_18__8_ (
		.chany_bottom_in(sb_1__1__297_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__298_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__345_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__345_chany_top_out[0:228]));

	cby_1__1_ cby_18__9_ (
		.chany_bottom_in(sb_1__1__298_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__299_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__346_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__346_chany_top_out[0:228]));

	cby_1__1_ cby_18__10_ (
		.chany_bottom_in(sb_1__1__299_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__300_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__347_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__347_chany_top_out[0:228]));

	cby_1__1_ cby_18__11_ (
		.chany_bottom_in(sb_1__1__300_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__301_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__348_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__348_chany_top_out[0:228]));

	cby_1__1_ cby_18__12_ (
		.chany_bottom_in(sb_1__1__301_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__302_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__349_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__349_chany_top_out[0:228]));

	cby_1__1_ cby_18__13_ (
		.chany_bottom_in(sb_1__1__302_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__303_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__350_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__350_chany_top_out[0:228]));

	cby_1__1_ cby_18__14_ (
		.chany_bottom_in(sb_1__1__303_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__304_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__351_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__351_chany_top_out[0:228]));

	cby_1__1_ cby_18__15_ (
		.chany_bottom_in(sb_1__1__304_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__305_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__352_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__352_chany_top_out[0:228]));

	cby_1__1_ cby_18__16_ (
		.chany_bottom_in(sb_1__1__305_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__306_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__353_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__353_chany_top_out[0:228]));

	cby_1__1_ cby_18__17_ (
		.chany_bottom_in(sb_1__1__306_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__307_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__354_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__354_chany_top_out[0:228]));

	cby_1__1_ cby_18__18_ (
		.chany_bottom_in(sb_1__1__307_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__308_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__355_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__355_chany_top_out[0:228]));

	cby_1__1_ cby_18__19_ (
		.chany_bottom_in(sb_1__1__308_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__309_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__356_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__356_chany_top_out[0:228]));

	cby_1__1_ cby_18__20_ (
		.chany_bottom_in(sb_1__1__309_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__310_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__357_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__357_chany_top_out[0:228]));

	cby_1__1_ cby_18__21_ (
		.chany_bottom_in(sb_1__1__310_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__311_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__358_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__358_chany_top_out[0:228]));

	cby_1__1_ cby_18__22_ (
		.chany_bottom_in(sb_1__1__311_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__17_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__359_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__359_chany_top_out[0:228]));

	cby_1__1_ cby_19__1_ (
		.chany_bottom_in(sb_1__0__18_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__312_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__360_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__360_chany_top_out[0:228]));

	cby_1__1_ cby_19__2_ (
		.chany_bottom_in(sb_1__1__312_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__313_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__361_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__361_chany_top_out[0:228]));

	cby_1__1_ cby_19__3_ (
		.chany_bottom_in(sb_1__1__313_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__314_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__362_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__362_chany_top_out[0:228]));

	cby_1__1_ cby_19__4_ (
		.chany_bottom_in(sb_1__1__314_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__18_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__363_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__363_chany_top_out[0:228]));

	cby_1__1_ cby_19__6_ (
		.chany_bottom_in(sb_1__5__12_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__315_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__364_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__364_chany_top_out[0:228]));

	cby_1__1_ cby_19__7_ (
		.chany_bottom_in(sb_1__1__315_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__316_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__365_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__365_chany_top_out[0:228]));

	cby_1__1_ cby_19__8_ (
		.chany_bottom_in(sb_1__1__316_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__317_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__366_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__366_chany_top_out[0:228]));

	cby_1__1_ cby_19__9_ (
		.chany_bottom_in(sb_1__1__317_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__318_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__367_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__367_chany_top_out[0:228]));

	cby_1__1_ cby_19__10_ (
		.chany_bottom_in(sb_1__1__318_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__319_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__368_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__368_chany_top_out[0:228]));

	cby_1__1_ cby_19__11_ (
		.chany_bottom_in(sb_1__1__319_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__320_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__369_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__369_chany_top_out[0:228]));

	cby_1__1_ cby_19__12_ (
		.chany_bottom_in(sb_1__1__320_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__321_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__370_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__370_chany_top_out[0:228]));

	cby_1__1_ cby_19__13_ (
		.chany_bottom_in(sb_1__1__321_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__322_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__371_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__371_chany_top_out[0:228]));

	cby_1__1_ cby_19__14_ (
		.chany_bottom_in(sb_1__1__322_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__323_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__372_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__372_chany_top_out[0:228]));

	cby_1__1_ cby_19__15_ (
		.chany_bottom_in(sb_1__1__323_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__324_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__373_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__373_chany_top_out[0:228]));

	cby_1__1_ cby_19__16_ (
		.chany_bottom_in(sb_1__1__324_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__325_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__374_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__374_chany_top_out[0:228]));

	cby_1__1_ cby_19__17_ (
		.chany_bottom_in(sb_1__1__325_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__326_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__375_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__375_chany_top_out[0:228]));

	cby_1__1_ cby_19__18_ (
		.chany_bottom_in(sb_1__1__326_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__327_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__376_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__376_chany_top_out[0:228]));

	cby_1__1_ cby_19__19_ (
		.chany_bottom_in(sb_1__1__327_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__328_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__377_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__377_chany_top_out[0:228]));

	cby_1__1_ cby_19__20_ (
		.chany_bottom_in(sb_1__1__328_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__329_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__378_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__378_chany_top_out[0:228]));

	cby_1__1_ cby_19__21_ (
		.chany_bottom_in(sb_1__1__329_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__330_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__379_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__379_chany_top_out[0:228]));

	cby_1__1_ cby_19__22_ (
		.chany_bottom_in(sb_1__1__330_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__18_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__380_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__380_chany_top_out[0:228]));

	cby_1__1_ cby_20__1_ (
		.chany_bottom_in(sb_1__0__19_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__331_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__381_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__381_chany_top_out[0:228]));

	cby_1__1_ cby_20__2_ (
		.chany_bottom_in(sb_1__1__331_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__332_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__382_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__382_chany_top_out[0:228]));

	cby_1__1_ cby_20__3_ (
		.chany_bottom_in(sb_1__1__332_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__333_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__383_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__383_chany_top_out[0:228]));

	cby_1__1_ cby_20__4_ (
		.chany_bottom_in(sb_1__1__333_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__19_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__384_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__384_chany_top_out[0:228]));

	cby_1__1_ cby_20__6_ (
		.chany_bottom_in(sb_1__5__13_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__334_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__385_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__385_chany_top_out[0:228]));

	cby_1__1_ cby_20__7_ (
		.chany_bottom_in(sb_1__1__334_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__335_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__386_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__386_chany_top_out[0:228]));

	cby_1__1_ cby_20__8_ (
		.chany_bottom_in(sb_1__1__335_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__336_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__387_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__387_chany_top_out[0:228]));

	cby_1__1_ cby_20__9_ (
		.chany_bottom_in(sb_1__1__336_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__337_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__388_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__388_chany_top_out[0:228]));

	cby_1__1_ cby_20__10_ (
		.chany_bottom_in(sb_1__1__337_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__338_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__389_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__389_chany_top_out[0:228]));

	cby_1__1_ cby_20__11_ (
		.chany_bottom_in(sb_1__1__338_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__339_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__390_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__390_chany_top_out[0:228]));

	cby_1__1_ cby_20__12_ (
		.chany_bottom_in(sb_1__1__339_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__340_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__391_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__391_chany_top_out[0:228]));

	cby_1__1_ cby_20__13_ (
		.chany_bottom_in(sb_1__1__340_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__341_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__392_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__392_chany_top_out[0:228]));

	cby_1__1_ cby_20__14_ (
		.chany_bottom_in(sb_1__1__341_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__342_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__393_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__393_chany_top_out[0:228]));

	cby_1__1_ cby_20__15_ (
		.chany_bottom_in(sb_1__1__342_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__343_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__394_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__394_chany_top_out[0:228]));

	cby_1__1_ cby_20__16_ (
		.chany_bottom_in(sb_1__1__343_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__344_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__395_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__395_chany_top_out[0:228]));

	cby_1__1_ cby_20__17_ (
		.chany_bottom_in(sb_1__1__344_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__345_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__396_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__396_chany_top_out[0:228]));

	cby_1__1_ cby_20__18_ (
		.chany_bottom_in(sb_1__1__345_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__346_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__397_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__397_chany_top_out[0:228]));

	cby_1__1_ cby_20__19_ (
		.chany_bottom_in(sb_1__1__346_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__347_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__398_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__398_chany_top_out[0:228]));

	cby_1__1_ cby_20__20_ (
		.chany_bottom_in(sb_1__1__347_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__348_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__399_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__399_chany_top_out[0:228]));

	cby_1__1_ cby_20__21_ (
		.chany_bottom_in(sb_1__1__348_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__349_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__400_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__400_chany_top_out[0:228]));

	cby_1__1_ cby_20__22_ (
		.chany_bottom_in(sb_1__1__349_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__19_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__401_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__401_chany_top_out[0:228]));

	cby_1__1_ cby_21__1_ (
		.chany_bottom_in(sb_1__0__20_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__350_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__402_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__402_chany_top_out[0:228]));

	cby_1__1_ cby_21__2_ (
		.chany_bottom_in(sb_1__1__350_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__351_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__403_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__403_chany_top_out[0:228]));

	cby_1__1_ cby_21__3_ (
		.chany_bottom_in(sb_1__1__351_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__352_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__404_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__404_chany_top_out[0:228]));

	cby_1__1_ cby_21__4_ (
		.chany_bottom_in(sb_1__1__352_chany_top_out[0:228]),
		.chany_top_in(sb_1__4__20_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__405_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__405_chany_top_out[0:228]));

	cby_1__1_ cby_21__6_ (
		.chany_bottom_in(sb_1__5__14_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__353_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__406_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__406_chany_top_out[0:228]));

	cby_1__1_ cby_21__7_ (
		.chany_bottom_in(sb_1__1__353_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__354_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__407_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__407_chany_top_out[0:228]));

	cby_1__1_ cby_21__8_ (
		.chany_bottom_in(sb_1__1__354_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__355_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__408_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__408_chany_top_out[0:228]));

	cby_1__1_ cby_21__9_ (
		.chany_bottom_in(sb_1__1__355_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__356_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__409_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__409_chany_top_out[0:228]));

	cby_1__1_ cby_21__10_ (
		.chany_bottom_in(sb_1__1__356_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__357_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__410_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__410_chany_top_out[0:228]));

	cby_1__1_ cby_21__11_ (
		.chany_bottom_in(sb_1__1__357_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__358_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__411_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__411_chany_top_out[0:228]));

	cby_1__1_ cby_21__12_ (
		.chany_bottom_in(sb_1__1__358_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__359_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__412_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__412_chany_top_out[0:228]));

	cby_1__1_ cby_21__13_ (
		.chany_bottom_in(sb_1__1__359_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__360_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__413_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__413_chany_top_out[0:228]));

	cby_1__1_ cby_21__14_ (
		.chany_bottom_in(sb_1__1__360_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__361_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__414_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__414_chany_top_out[0:228]));

	cby_1__1_ cby_21__15_ (
		.chany_bottom_in(sb_1__1__361_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__362_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__415_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__415_chany_top_out[0:228]));

	cby_1__1_ cby_21__16_ (
		.chany_bottom_in(sb_1__1__362_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__363_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__416_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__416_chany_top_out[0:228]));

	cby_1__1_ cby_21__17_ (
		.chany_bottom_in(sb_1__1__363_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__364_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__417_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__417_chany_top_out[0:228]));

	cby_1__1_ cby_21__18_ (
		.chany_bottom_in(sb_1__1__364_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__365_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__418_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__418_chany_top_out[0:228]));

	cby_1__1_ cby_21__19_ (
		.chany_bottom_in(sb_1__1__365_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__366_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__419_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__419_chany_top_out[0:228]));

	cby_1__1_ cby_21__20_ (
		.chany_bottom_in(sb_1__1__366_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__367_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__420_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__420_chany_top_out[0:228]));

	cby_1__1_ cby_21__21_ (
		.chany_bottom_in(sb_1__1__367_chany_top_out[0:228]),
		.chany_top_in(sb_1__1__368_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__421_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__421_chany_top_out[0:228]));

	cby_1__1_ cby_21__22_ (
		.chany_bottom_in(sb_1__1__368_chany_top_out[0:228]),
		.chany_top_in(sb_1__22__20_chany_bottom_out[0:228]),
		.chany_bottom_out(cby_1__1__422_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__1__422_chany_top_out[0:228]));

	cby_1__5_ cby_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__0_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__0_ccff_tail),
		.chany_bottom_out(cby_1__5__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__0_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__0_ccff_tail));

	cby_1__5_ cby_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__1_chany_top_out[0:228]),
		.chany_top_in(sb_2__5__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__1_ccff_tail),
		.chany_bottom_out(cby_1__5__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__1_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__1_ccff_tail));

	cby_1__5_ cby_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__2_chany_top_out[0:228]),
		.chany_top_in(sb_3__5__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__2_ccff_tail),
		.chany_bottom_out(cby_1__5__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__2_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__2_ccff_tail));

	cby_1__5_ cby_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__3_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__1_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__3_ccff_tail),
		.chany_bottom_out(cby_1__5__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__3_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__3_ccff_tail));

	cby_1__5_ cby_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__4_chany_top_out[0:228]),
		.chany_top_in(sb_2__5__1_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__4_ccff_tail),
		.chany_bottom_out(cby_1__5__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__4_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__4_ccff_tail));

	cby_1__5_ cby_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__5_chany_top_out[0:228]),
		.chany_top_in(sb_3__5__1_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__5_ccff_tail),
		.chany_bottom_out(cby_1__5__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__5_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__5_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__5_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__5_ccff_tail));

	cby_1__5_ cby_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__6_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__2_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__6_ccff_tail),
		.chany_bottom_out(cby_1__5__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__6_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__6_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__6_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__6_ccff_tail));

	cby_1__5_ cby_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__7_chany_top_out[0:228]),
		.chany_top_in(sb_2__5__2_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__7_ccff_tail),
		.chany_bottom_out(cby_1__5__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__7_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__7_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__7_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__7_ccff_tail));

	cby_1__5_ cby_9__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__8_chany_top_out[0:228]),
		.chany_top_in(sb_3__5__2_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__8_ccff_tail),
		.chany_bottom_out(cby_1__5__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__8_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__8_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__8_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__8_ccff_tail));

	cby_1__5_ cby_10__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__9_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__3_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__9_ccff_tail),
		.chany_bottom_out(cby_1__5__9_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__9_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__9_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__9_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__9_ccff_tail));

	cby_1__5_ cby_11__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__10_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__4_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__10_ccff_tail),
		.chany_bottom_out(cby_1__5__10_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__10_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__10_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__10_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__10_ccff_tail));

	cby_1__5_ cby_12__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__11_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__5_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__11_ccff_tail),
		.chany_bottom_out(cby_1__5__11_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__11_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__11_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__11_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__11_ccff_tail));

	cby_1__5_ cby_13__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__12_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__6_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__12_ccff_tail),
		.chany_bottom_out(cby_1__5__12_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__12_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__12_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__12_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__12_ccff_tail));

	cby_1__5_ cby_14__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__13_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__7_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__13_ccff_tail),
		.chany_bottom_out(cby_1__5__13_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__13_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__13_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__13_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__13_ccff_tail));

	cby_1__5_ cby_15__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__14_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__8_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__14_ccff_tail),
		.chany_bottom_out(cby_1__5__14_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__14_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__14_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__14_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__14_ccff_tail));

	cby_1__5_ cby_16__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__15_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__9_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__15_ccff_tail),
		.chany_bottom_out(cby_1__5__15_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__15_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__15_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__15_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__15_ccff_tail));

	cby_1__5_ cby_17__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__16_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__10_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__16_ccff_tail),
		.chany_bottom_out(cby_1__5__16_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__16_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__16_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__16_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__16_ccff_tail));

	cby_1__5_ cby_18__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__17_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__11_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__17_ccff_tail),
		.chany_bottom_out(cby_1__5__17_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__17_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__17_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__17_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__17_ccff_tail));

	cby_1__5_ cby_19__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__18_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__12_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__18_ccff_tail),
		.chany_bottom_out(cby_1__5__18_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__18_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__18_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__18_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__18_ccff_tail));

	cby_1__5_ cby_20__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__19_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__13_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__19_ccff_tail),
		.chany_bottom_out(cby_1__5__19_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__19_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__19_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__19_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__19_ccff_tail));

	cby_1__5_ cby_21__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__4__20_chany_top_out[0:228]),
		.chany_top_in(sb_1__5__14_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__20_ccff_tail),
		.chany_bottom_out(cby_1__5__20_chany_bottom_out[0:228]),
		.chany_top_out(cby_1__5__20_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__5__20_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__5__20_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__5__20_ccff_tail));

	cby_2__3_ cby_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__0_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__0_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__0_ccff_tail),
		.chany_bottom_out(cby_2__3__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__0_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__0_ccff_tail));

	cby_2__3_ cby_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__5__0_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__1_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__5__1_ccff_tail),
		.chany_bottom_out(cby_2__3__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__1_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__1_ccff_tail));

	cby_2__3_ cby_2__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__1_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__2_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__1_ccff_tail),
		.chany_bottom_out(cby_2__3__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__2_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__2_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__2_ccff_tail));

	cby_2__3_ cby_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__2_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__3_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__2_ccff_tail),
		.chany_bottom_out(cby_2__3__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__3_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__3_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__3_ccff_tail));

	cby_2__3_ cby_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__5__1_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__4_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__5__3_ccff_tail),
		.chany_bottom_out(cby_2__3__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__4_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__4_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__4_ccff_tail));

	cby_2__3_ cby_5__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__3_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__5_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__3_ccff_tail),
		.chany_bottom_out(cby_2__3__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__5_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__5_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__5_ccff_tail));

	cby_2__3_ cby_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__4_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__6_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__4_ccff_tail),
		.chany_bottom_out(cby_2__3__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__6_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__6_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__6_ccff_tail));

	cby_2__3_ cby_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__5__2_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__7_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__5__5_ccff_tail),
		.chany_bottom_out(cby_2__3__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__7_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__7_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__7_ccff_tail));

	cby_2__3_ cby_8__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__2__5_chany_top_out[0:228]),
		.chany_top_in(sb_2__3__8_chany_bottom_out[0:228]),
		.ccff_head(sb_2__2__5_ccff_tail),
		.chany_bottom_out(cby_2__3__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_2__3__8_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_2__3__8_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.ccff_tail(cby_2__3__8_ccff_tail));

	cby_3__3_ cby_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__0_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__0_ccff_tail),
		.chany_bottom_out(cby_3__3__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__0_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__0_ccff_tail));

	cby_3__3_ cby_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__5__0_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__1_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__5__0_ccff_tail),
		.chany_bottom_out(cby_3__3__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__1_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__1_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__1_ccff_tail));

	cby_3__3_ cby_3__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__1_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__2_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__1_ccff_tail),
		.chany_bottom_out(cby_3__3__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__2_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__2_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__2_ccff_tail));

	cby_3__3_ cby_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__2_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__3_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__2_ccff_tail),
		.chany_bottom_out(cby_3__3__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__3_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__3_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__3_ccff_tail));

	cby_3__3_ cby_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__5__1_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__4_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__5__1_ccff_tail),
		.chany_bottom_out(cby_3__3__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__4_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__4_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__4_ccff_tail));

	cby_3__3_ cby_6__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__3_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__5_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__3_ccff_tail),
		.chany_bottom_out(cby_3__3__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__5_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__5_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__5_ccff_tail));

	cby_3__3_ cby_9__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__4_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__6_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__4_ccff_tail),
		.chany_bottom_out(cby_3__3__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__6_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__6_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__6_ccff_tail));

	cby_3__3_ cby_9__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__5__2_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__7_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__5__2_ccff_tail),
		.chany_bottom_out(cby_3__3__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__7_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__7_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__7_ccff_tail));

	cby_3__3_ cby_9__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__5_chany_top_out[0:228]),
		.chany_top_in(sb_3__3__8_chany_bottom_out[0:228]),
		.ccff_head(cbx_3__2__5_ccff_tail),
		.chany_bottom_out(cby_3__3__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_3__3__8_chany_top_out[0:228]),
		.left_grid_right_width_0_height_0_subtile_0__pin_rst__0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_rst__0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_3__3__8_left_grid_right_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.ccff_tail(cby_3__3__8_ccff_tail));

	cby_22__1_ cby_22__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__0__0_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__0__21_ccff_tail),
		.chany_bottom_out(cby_22__1__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__0_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__0_ccff_tail));

	cby_22__1_ cby_22__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__0_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__1_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__0_ccff_tail),
		.chany_bottom_out(cby_22__1__1_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__1_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__1_ccff_tail));

	cby_22__1_ cby_22__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__1_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__2_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__1_ccff_tail),
		.chany_bottom_out(cby_22__1__2_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__2_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__2_ccff_tail));

	cby_22__1_ cby_22__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__2_chany_top_out[0:228]),
		.chany_top_in(sb_22__4__0_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__2_ccff_tail),
		.chany_bottom_out(cby_22__1__3_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__3_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__3_ccff_tail));

	cby_22__1_ cby_22__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__5__0_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__3_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__5__18_ccff_tail),
		.chany_bottom_out(cby_22__1__4_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__4_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__4_ccff_tail));

	cby_22__1_ cby_22__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__3_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__4_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__3_ccff_tail),
		.chany_bottom_out(cby_22__1__5_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__5_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__5_ccff_tail));

	cby_22__1_ cby_22__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__4_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__5_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__4_ccff_tail),
		.chany_bottom_out(cby_22__1__6_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__6_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__6_ccff_tail));

	cby_22__1_ cby_22__9_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__5_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__6_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__5_ccff_tail),
		.chany_bottom_out(cby_22__1__7_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__7_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__7_ccff_tail));

	cby_22__1_ cby_22__10_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__6_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__7_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__6_ccff_tail),
		.chany_bottom_out(cby_22__1__8_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__8_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__8_ccff_tail));

	cby_22__1_ cby_22__11_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__7_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__8_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__7_ccff_tail),
		.chany_bottom_out(cby_22__1__9_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__9_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__9_ccff_tail));

	cby_22__1_ cby_22__12_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__8_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__9_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__8_ccff_tail),
		.chany_bottom_out(cby_22__1__10_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__10_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__10_ccff_tail));

	cby_22__1_ cby_22__13_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__9_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__10_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__9_ccff_tail),
		.chany_bottom_out(cby_22__1__11_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__11_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__11_ccff_tail));

	cby_22__1_ cby_22__14_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__10_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__11_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__10_ccff_tail),
		.chany_bottom_out(cby_22__1__12_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__12_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__12_ccff_tail));

	cby_22__1_ cby_22__15_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__11_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__12_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__11_ccff_tail),
		.chany_bottom_out(cby_22__1__13_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__13_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__13_ccff_tail));

	cby_22__1_ cby_22__16_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__12_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__13_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__12_ccff_tail),
		.chany_bottom_out(cby_22__1__14_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__14_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__14_ccff_tail));

	cby_22__1_ cby_22__17_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__13_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__14_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__13_ccff_tail),
		.chany_bottom_out(cby_22__1__15_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__15_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__15_ccff_tail));

	cby_22__1_ cby_22__18_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__14_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__15_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__14_ccff_tail),
		.chany_bottom_out(cby_22__1__16_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__16_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__16_ccff_tail));

	cby_22__1_ cby_22__19_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__15_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__16_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__15_ccff_tail),
		.chany_bottom_out(cby_22__1__17_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__17_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__17_ccff_tail));

	cby_22__1_ cby_22__20_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__16_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__17_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__16_ccff_tail),
		.chany_bottom_out(cby_22__1__18_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__18_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__18_ccff_tail));

	cby_22__1_ cby_22__21_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__17_chany_top_out[0:228]),
		.chany_top_in(sb_22__1__18_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__17_ccff_tail),
		.chany_bottom_out(cby_22__1__19_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__19_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__19_ccff_tail));

	cby_22__1_ cby_22__22_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__1__18_chany_top_out[0:228]),
		.chany_top_in(sb_22__22__0_chany_bottom_out[0:228]),
		.ccff_head(sb_22__1__18_ccff_tail),
		.chany_bottom_out(cby_22__1__20_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__1__20_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_22__1__20_ccff_tail));

	cby_22__5_ cby_22__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_22__4__0_chany_top_out[0:228]),
		.chany_top_in(sb_22__5__0_chany_bottom_out[0:228]),
		.ccff_head(cbx_1__4__21_ccff_tail),
		.chany_bottom_out(cby_22__5__0_chany_bottom_out[0:228]),
		.chany_top_out(cby_22__5__0_chany_top_out[0:228]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_22__5__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_22__5__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_22__5__0_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




