//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[3][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Sep  9 09:18:43 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_3__2_ -----
module sb_3__2_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_,
                chanx_right_in,
                chany_bottom_in,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:166] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_;
//----- INPUT PORTS -----
input [0:166] chanx_right_in;
//----- INPUT PORTS -----
input [0:166] chany_bottom_in;
//----- INPUT PORTS -----
input [0:166] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:166] chany_top_out;
//----- OUTPUT PORTS -----
output [0:166] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:166] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:166] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size13_0_sram;
wire [0:7] mux_2level_tapbuf_size13_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_1_sram;
wire [0:7] mux_2level_tapbuf_size13_1_sram_inv;
wire [0:0] mux_2level_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_1_ccff_tail;
wire [0:7] mux_2level_tapbuf_size14_0_sram;
wire [0:7] mux_2level_tapbuf_size14_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_10_sram;
wire [0:7] mux_2level_tapbuf_size14_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_11_sram;
wire [0:7] mux_2level_tapbuf_size14_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_12_sram;
wire [0:7] mux_2level_tapbuf_size14_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_13_sram;
wire [0:7] mux_2level_tapbuf_size14_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_14_sram;
wire [0:7] mux_2level_tapbuf_size14_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_15_sram;
wire [0:7] mux_2level_tapbuf_size14_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_16_sram;
wire [0:7] mux_2level_tapbuf_size14_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_17_sram;
wire [0:7] mux_2level_tapbuf_size14_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_18_sram;
wire [0:7] mux_2level_tapbuf_size14_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_19_sram;
wire [0:7] mux_2level_tapbuf_size14_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_1_sram;
wire [0:7] mux_2level_tapbuf_size14_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_20_sram;
wire [0:7] mux_2level_tapbuf_size14_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_21_sram;
wire [0:7] mux_2level_tapbuf_size14_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_22_sram;
wire [0:7] mux_2level_tapbuf_size14_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_23_sram;
wire [0:7] mux_2level_tapbuf_size14_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_24_sram;
wire [0:7] mux_2level_tapbuf_size14_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_25_sram;
wire [0:7] mux_2level_tapbuf_size14_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_26_sram;
wire [0:7] mux_2level_tapbuf_size14_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_27_sram;
wire [0:7] mux_2level_tapbuf_size14_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_28_sram;
wire [0:7] mux_2level_tapbuf_size14_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_29_sram;
wire [0:7] mux_2level_tapbuf_size14_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_2_sram;
wire [0:7] mux_2level_tapbuf_size14_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_30_sram;
wire [0:7] mux_2level_tapbuf_size14_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_31_sram;
wire [0:7] mux_2level_tapbuf_size14_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_32_sram;
wire [0:7] mux_2level_tapbuf_size14_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_33_sram;
wire [0:7] mux_2level_tapbuf_size14_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_34_sram;
wire [0:7] mux_2level_tapbuf_size14_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_35_sram;
wire [0:7] mux_2level_tapbuf_size14_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_36_sram;
wire [0:7] mux_2level_tapbuf_size14_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_37_sram;
wire [0:7] mux_2level_tapbuf_size14_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_38_sram;
wire [0:7] mux_2level_tapbuf_size14_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_39_sram;
wire [0:7] mux_2level_tapbuf_size14_39_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_3_sram;
wire [0:7] mux_2level_tapbuf_size14_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_40_sram;
wire [0:7] mux_2level_tapbuf_size14_40_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_41_sram;
wire [0:7] mux_2level_tapbuf_size14_41_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_42_sram;
wire [0:7] mux_2level_tapbuf_size14_42_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_43_sram;
wire [0:7] mux_2level_tapbuf_size14_43_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_44_sram;
wire [0:7] mux_2level_tapbuf_size14_44_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_45_sram;
wire [0:7] mux_2level_tapbuf_size14_45_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_46_sram;
wire [0:7] mux_2level_tapbuf_size14_46_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_47_sram;
wire [0:7] mux_2level_tapbuf_size14_47_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_48_sram;
wire [0:7] mux_2level_tapbuf_size14_48_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_49_sram;
wire [0:7] mux_2level_tapbuf_size14_49_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_4_sram;
wire [0:7] mux_2level_tapbuf_size14_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_50_sram;
wire [0:7] mux_2level_tapbuf_size14_50_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_51_sram;
wire [0:7] mux_2level_tapbuf_size14_51_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_52_sram;
wire [0:7] mux_2level_tapbuf_size14_52_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_53_sram;
wire [0:7] mux_2level_tapbuf_size14_53_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_54_sram;
wire [0:7] mux_2level_tapbuf_size14_54_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_55_sram;
wire [0:7] mux_2level_tapbuf_size14_55_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_56_sram;
wire [0:7] mux_2level_tapbuf_size14_56_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_57_sram;
wire [0:7] mux_2level_tapbuf_size14_57_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_58_sram;
wire [0:7] mux_2level_tapbuf_size14_58_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_59_sram;
wire [0:7] mux_2level_tapbuf_size14_59_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_5_sram;
wire [0:7] mux_2level_tapbuf_size14_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_60_sram;
wire [0:7] mux_2level_tapbuf_size14_60_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_61_sram;
wire [0:7] mux_2level_tapbuf_size14_61_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_62_sram;
wire [0:7] mux_2level_tapbuf_size14_62_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_63_sram;
wire [0:7] mux_2level_tapbuf_size14_63_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_64_sram;
wire [0:7] mux_2level_tapbuf_size14_64_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_65_sram;
wire [0:7] mux_2level_tapbuf_size14_65_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_66_sram;
wire [0:7] mux_2level_tapbuf_size14_66_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_67_sram;
wire [0:7] mux_2level_tapbuf_size14_67_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_68_sram;
wire [0:7] mux_2level_tapbuf_size14_68_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_69_sram;
wire [0:7] mux_2level_tapbuf_size14_69_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_6_sram;
wire [0:7] mux_2level_tapbuf_size14_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_70_sram;
wire [0:7] mux_2level_tapbuf_size14_70_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_71_sram;
wire [0:7] mux_2level_tapbuf_size14_71_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_7_sram;
wire [0:7] mux_2level_tapbuf_size14_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_8_sram;
wire [0:7] mux_2level_tapbuf_size14_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size14_9_sram;
wire [0:7] mux_2level_tapbuf_size14_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size14_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size14_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size15_0_sram;
wire [0:7] mux_2level_tapbuf_size15_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_1_sram;
wire [0:7] mux_2level_tapbuf_size15_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_2_sram;
wire [0:7] mux_2level_tapbuf_size15_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_3_sram;
wire [0:7] mux_2level_tapbuf_size15_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_4_sram;
wire [0:7] mux_2level_tapbuf_size15_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_5_sram;
wire [0:7] mux_2level_tapbuf_size15_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_6_sram;
wire [0:7] mux_2level_tapbuf_size15_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_7_sram;
wire [0:7] mux_2level_tapbuf_size15_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_8_sram;
wire [0:7] mux_2level_tapbuf_size15_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size15_9_sram;
wire [0:7] mux_2level_tapbuf_size15_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size15_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_16_sram;
wire [0:5] mux_2level_tapbuf_size8_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_17_sram;
wire [0:5] mux_2level_tapbuf_size8_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_18_sram;
wire [0:5] mux_2level_tapbuf_size8_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_19_sram;
wire [0:5] mux_2level_tapbuf_size8_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_20_sram;
wire [0:5] mux_2level_tapbuf_size8_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_21_sram;
wire [0:5] mux_2level_tapbuf_size8_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_22_sram;
wire [0:5] mux_2level_tapbuf_size8_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_23_sram;
wire [0:5] mux_2level_tapbuf_size8_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_24_sram;
wire [0:5] mux_2level_tapbuf_size8_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_25_sram;
wire [0:5] mux_2level_tapbuf_size8_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_26_sram;
wire [0:5] mux_2level_tapbuf_size8_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_27_sram;
wire [0:5] mux_2level_tapbuf_size8_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_28_sram;
wire [0:5] mux_2level_tapbuf_size8_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_29_sram;
wire [0:5] mux_2level_tapbuf_size8_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_30_sram;
wire [0:5] mux_2level_tapbuf_size8_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_31_sram;
wire [0:5] mux_2level_tapbuf_size8_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_32_sram;
wire [0:5] mux_2level_tapbuf_size8_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_33_sram;
wire [0:5] mux_2level_tapbuf_size8_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_34_sram;
wire [0:5] mux_2level_tapbuf_size8_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_35_sram;
wire [0:5] mux_2level_tapbuf_size8_35_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_36_sram;
wire [0:5] mux_2level_tapbuf_size8_36_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_37_sram;
wire [0:5] mux_2level_tapbuf_size8_37_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_38_sram;
wire [0:5] mux_2level_tapbuf_size8_38_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_39_sram;
wire [0:5] mux_2level_tapbuf_size8_39_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_40_sram;
wire [0:5] mux_2level_tapbuf_size8_40_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_41_sram;
wire [0:5] mux_2level_tapbuf_size8_41_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_42_sram;
wire [0:5] mux_2level_tapbuf_size8_42_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_43_sram;
wire [0:5] mux_2level_tapbuf_size8_43_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_44_sram;
wire [0:5] mux_2level_tapbuf_size8_44_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_45_sram;
wire [0:5] mux_2level_tapbuf_size8_45_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_46_sram;
wire [0:5] mux_2level_tapbuf_size8_46_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_47_sram;
wire [0:5] mux_2level_tapbuf_size8_47_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_48_sram;
wire [0:5] mux_2level_tapbuf_size8_48_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_49_sram;
wire [0:5] mux_2level_tapbuf_size8_49_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_50_sram;
wire [0:5] mux_2level_tapbuf_size8_50_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_51_sram;
wire [0:5] mux_2level_tapbuf_size8_51_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_52_sram;
wire [0:5] mux_2level_tapbuf_size8_52_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_53_sram;
wire [0:5] mux_2level_tapbuf_size8_53_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_54_sram;
wire [0:5] mux_2level_tapbuf_size8_54_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_55_sram;
wire [0:5] mux_2level_tapbuf_size8_55_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_56_sram;
wire [0:5] mux_2level_tapbuf_size8_56_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_57_sram;
wire [0:5] mux_2level_tapbuf_size8_57_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_58_sram;
wire [0:5] mux_2level_tapbuf_size8_58_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_59_sram;
wire [0:5] mux_2level_tapbuf_size8_59_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_60_sram;
wire [0:5] mux_2level_tapbuf_size8_60_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_61_sram;
wire [0:5] mux_2level_tapbuf_size8_61_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_62_sram;
wire [0:5] mux_2level_tapbuf_size8_62_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_63_sram;
wire [0:5] mux_2level_tapbuf_size8_63_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_64_sram;
wire [0:5] mux_2level_tapbuf_size8_64_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_65_sram;
wire [0:5] mux_2level_tapbuf_size8_65_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_66_sram;
wire [0:5] mux_2level_tapbuf_size8_66_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_67_sram;
wire [0:5] mux_2level_tapbuf_size8_67_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_68_sram;
wire [0:5] mux_2level_tapbuf_size8_68_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_69_sram;
wire [0:5] mux_2level_tapbuf_size8_69_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_70_sram;
wire [0:5] mux_2level_tapbuf_size8_70_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_71_sram;
wire [0:5] mux_2level_tapbuf_size8_71_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_72_sram;
wire [0:5] mux_2level_tapbuf_size8_72_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_73_sram;
wire [0:5] mux_2level_tapbuf_size8_73_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_74_sram;
wire [0:5] mux_2level_tapbuf_size8_74_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_75_sram;
wire [0:5] mux_2level_tapbuf_size8_75_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_76_sram;
wire [0:5] mux_2level_tapbuf_size8_76_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_77_sram;
wire [0:5] mux_2level_tapbuf_size8_77_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_78_sram;
wire [0:5] mux_2level_tapbuf_size8_78_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_79_sram;
wire [0:5] mux_2level_tapbuf_size8_79_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size15 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[57], chanx_right_in[113], chanx_left_in[0], chanx_left_in[3], chanx_left_in[56], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size15_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_0_sram_inv[0:7]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size15 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[12], chanx_right_in[39], chanx_right_in[68], chanx_right_in[124], chanx_left_in[45], chanx_left_in[101], chanx_left_in[139], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size15_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_1_sram_inv[0:7]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size15 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[22], chanx_right_in[71], chanx_right_in[78], chanx_right_in[134], chanx_left_in[34], chanx_left_in[90], chanx_left_in[107], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size15_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_2_sram_inv[0:7]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size15 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[33], chanx_right_in[89], chanx_right_in[103], chanx_right_in[145], chanx_left_in[24], chanx_left_in[75], chanx_left_in[80], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size15_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_3_sram_inv[0:7]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size15 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[44], chanx_right_in[100], chanx_right_in[135], chanx_right_in[156], chanx_left_in[13], chanx_left_in[43], chanx_left_in[69], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size15_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_4_sram_inv[0:7]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size15 mux_left_track_65 (
		.in({chany_top_in[45], chany_top_in[101], chany_top_in[139], chany_top_in[157], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[65], chany_bottom_in[121], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size15_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_5_sram_inv[0:7]),
		.out(chanx_left_out[32]));

	mux_2level_tapbuf_size15 mux_left_track_129 (
		.in({chany_top_in[34], chany_top_in[90], chany_top_in[107], chany_top_in[146], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[76], chany_bottom_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size15_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_6_sram_inv[0:7]),
		.out(chanx_left_out[64]));

	mux_2level_tapbuf_size15 mux_left_track_193 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[80], chany_top_in[136], chany_bottom_in[30], chany_bottom_in[86], chany_bottom_in[95], chany_bottom_in[142], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size15_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_7_sram_inv[0:7]),
		.out(chanx_left_out[96]));

	mux_2level_tapbuf_size15 mux_left_track_257 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[69], chany_top_in[125], chany_bottom_in[41], chany_bottom_in[97], chany_bottom_in[127], chany_bottom_in[153], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size15_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_8_sram_inv[0:7]),
		.out(chanx_left_out[128]));

	mux_2level_tapbuf_size15 mux_left_track_321 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[58], chany_top_in[114], chany_bottom_in[52], chany_bottom_in[108], chany_bottom_in[159], chany_bottom_in[164], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size15_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_9_sram_inv[0:7]),
		.out(chanx_left_out[160]));

	mux_2level_tapbuf_size15_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_0_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_1_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_2_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_3_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_4_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_left_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_5_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_left_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_6_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_left_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_7_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_left_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_8_sram_inv[0:7]));

	mux_2level_tapbuf_size15_mem mem_left_track_321 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_9_sram_inv[0:7]));

	mux_2level_tapbuf_size13 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[58], chanx_right_in[114], chanx_left_in[54], chanx_left_in[110], chanx_left_in[166]}),
		.sram(mux_2level_tapbuf_size13_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_0_sram_inv[0:7]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size13 mux_left_track_9 (
		.in({chany_top_in[54], chany_top_in[110], chany_top_in[166], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[56], chany_bottom_in[112], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_}),
		.sram(mux_2level_tapbuf_size13_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_1_sram_inv[0:7]),
		.out(chanx_left_out[4]));

	mux_2level_tapbuf_size13_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_0_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_left_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_1_sram_inv[0:7]));

	mux_2level_tapbuf_size14 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[4], chanx_right_in[15], chanx_right_in[60], chanx_right_in[116], chanx_left_in[53], chanx_left_in[109], chanx_left_in[163], chanx_left_in[165]}),
		.sram(mux_2level_tapbuf_size14_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_0_sram_inv[0:7]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size14 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, chanx_right_in[5], chanx_right_in[19], chanx_right_in[61], chanx_right_in[117], chanx_left_in[52], chanx_left_in[108], chanx_left_in[159], chanx_left_in[164]}),
		.sram(mux_2level_tapbuf_size14_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_1_sram_inv[0:7]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size14 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, chanx_right_in[6], chanx_right_in[23], chanx_right_in[62], chanx_right_in[118], chanx_left_in[50], chanx_left_in[106], chanx_left_in[155], chanx_left_in[162]}),
		.sram(mux_2level_tapbuf_size14_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_2_sram_inv[0:7]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size14 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[64], chanx_right_in[120], chanx_left_in[49], chanx_left_in[105], chanx_left_in[151], chanx_left_in[161]}),
		.sram(mux_2level_tapbuf_size14_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_3_sram_inv[0:7]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size14 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_right_in[9], chanx_right_in[31], chanx_right_in[65], chanx_right_in[121], chanx_left_in[48], chanx_left_in[104], chanx_left_in[147], chanx_left_in[160]}),
		.sram(mux_2level_tapbuf_size14_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_4_sram_inv[0:7]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size14 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[10], chanx_right_in[35], chanx_right_in[66], chanx_right_in[122], chanx_left_in[46], chanx_left_in[102], chanx_left_in[143], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size14_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_5_sram_inv[0:7]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size14 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, chanx_right_in[13], chanx_right_in[43], chanx_right_in[69], chanx_right_in[125], chanx_left_in[44], chanx_left_in[100], chanx_left_in[135], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size14_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_6_sram_inv[0:7]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size14 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[14], chanx_right_in[47], chanx_right_in[70], chanx_right_in[126], chanx_left_in[42], chanx_left_in[98], chanx_left_in[131], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size14_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_7_sram_inv[0:7]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size14 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, chanx_right_in[16], chanx_right_in[51], chanx_right_in[72], chanx_right_in[128], chanx_left_in[41], chanx_left_in[97], chanx_left_in[127], chanx_left_in[153]}),
		.sram(mux_2level_tapbuf_size14_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_8_sram_inv[0:7]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size14 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, chanx_right_in[17], chanx_right_in[55], chanx_right_in[73], chanx_right_in[129], chanx_left_in[40], chanx_left_in[96], chanx_left_in[123], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size14_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_9_sram_inv[0:7]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size14 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[18], chanx_right_in[59], chanx_right_in[74], chanx_right_in[130], chanx_left_in[38], chanx_left_in[94], chanx_left_in[119], chanx_left_in[150]}),
		.sram(mux_2level_tapbuf_size14_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_10_sram_inv[0:7]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size14 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_right_in[20], chanx_right_in[63], chanx_right_in[76], chanx_right_in[132], chanx_left_in[37], chanx_left_in[93], chanx_left_in[115], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size14_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_11_sram_inv[0:7]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size14 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[21], chanx_right_in[67], chanx_right_in[77], chanx_right_in[133], chanx_left_in[36], chanx_left_in[92], chanx_left_in[111], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size14_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_12_sram_inv[0:7]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size14 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, chanx_right_in[24], chanx_right_in[75], chanx_right_in[80], chanx_right_in[136], chanx_left_in[33], chanx_left_in[89], chanx_left_in[103], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size14_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_13_sram_inv[0:7]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size14 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[25], chanx_right_in[79], chanx_right_in[81], chanx_right_in[137], chanx_left_in[32], chanx_left_in[88], chanx_left_in[99], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size14_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_14_sram_inv[0:7]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size14 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, chanx_right_in[26], chanx_right_in[82:83], chanx_right_in[138], chanx_left_in[30], chanx_left_in[86], chanx_left_in[95], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size14_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_15_sram_inv[0:7]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size14 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, chanx_right_in[28], chanx_right_in[84], chanx_right_in[87], chanx_right_in[140], chanx_left_in[29], chanx_left_in[85], chanx_left_in[91], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size14_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_16_sram_inv[0:7]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size14 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[29], chanx_right_in[85], chanx_right_in[91], chanx_right_in[141], chanx_left_in[28], chanx_left_in[84], chanx_left_in[87], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size14_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_17_sram_inv[0:7]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size14 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_right_in[30], chanx_right_in[86], chanx_right_in[95], chanx_right_in[142], chanx_left_in[26], chanx_left_in[82:83], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size14_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_18_sram_inv[0:7]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size14 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[32], chanx_right_in[88], chanx_right_in[99], chanx_right_in[144], chanx_left_in[25], chanx_left_in[79], chanx_left_in[81], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size14_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_19_sram_inv[0:7]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size14 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, chanx_right_in[34], chanx_right_in[90], chanx_right_in[107], chanx_right_in[146], chanx_left_in[22], chanx_left_in[71], chanx_left_in[78], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size14_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_20_sram_inv[0:7]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size14 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[36], chanx_right_in[92], chanx_right_in[111], chanx_right_in[148], chanx_left_in[21], chanx_left_in[67], chanx_left_in[77], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size14_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_21_sram_inv[0:7]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size14 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, chanx_right_in[37], chanx_right_in[93], chanx_right_in[115], chanx_right_in[149], chanx_left_in[20], chanx_left_in[63], chanx_left_in[76], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size14_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_22_sram_inv[0:7]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size14 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, chanx_right_in[38], chanx_right_in[94], chanx_right_in[119], chanx_right_in[150], chanx_left_in[18], chanx_left_in[59], chanx_left_in[74], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size14_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_23_sram_inv[0:7]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size14 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[40], chanx_right_in[96], chanx_right_in[123], chanx_right_in[152], chanx_left_in[17], chanx_left_in[55], chanx_left_in[73], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size14_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_24_sram_inv[0:7]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size14 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_right_in[41], chanx_right_in[97], chanx_right_in[127], chanx_right_in[153], chanx_left_in[16], chanx_left_in[51], chanx_left_in[72], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size14_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_25_sram_inv[0:7]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size14 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[42], chanx_right_in[98], chanx_right_in[131], chanx_right_in[154], chanx_left_in[14], chanx_left_in[47], chanx_left_in[70], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size14_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_26_sram_inv[0:7]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size14 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, chanx_right_in[45], chanx_right_in[101], chanx_right_in[139], chanx_right_in[157], chanx_left_in[12], chanx_left_in[39], chanx_left_in[68], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size14_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_27_sram_inv[0:7]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size14 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_18_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_26_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_34_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[46], chanx_right_in[102], chanx_right_in[143], chanx_right_in[158], chanx_left_in[10], chanx_left_in[35], chanx_left_in[66], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size14_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_28_sram_inv[0:7]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size14 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_19_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_27_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, chanx_right_in[48], chanx_right_in[104], chanx_right_in[147], chanx_right_in[160], chanx_left_in[9], chanx_left_in[31], chanx_left_in[65], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size14_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_29_sram_inv[0:7]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size14 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_, top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, chanx_right_in[49], chanx_right_in[105], chanx_right_in[151], chanx_right_in[161], chanx_left_in[8], chanx_left_in[27], chanx_left_in[64], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size14_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_30_sram_inv[0:7]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size14 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_21_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_29_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[50], chanx_right_in[106], chanx_right_in[155], chanx_right_in[162], chanx_left_in[6], chanx_left_in[23], chanx_left_in[62], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size14_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_31_sram_inv[0:7]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size14 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_14_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_22_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_30_, top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_right_in[52], chanx_right_in[108], chanx_right_in[159], chanx_right_in[164], chanx_left_in[5], chanx_left_in[19], chanx_left_in[61], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size14_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_32_sram_inv[0:7]),
		.out(chany_top_out[152]));

	mux_2level_tapbuf_size14 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_15_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_23_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_31_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[53], chanx_right_in[109], chanx_right_in[163], chanx_right_in[165], chanx_left_in[4], chanx_left_in[15], chanx_left_in[60], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size14_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_33_sram_inv[0:7]),
		.out(chany_top_out[156]));

	mux_2level_tapbuf_size14 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_, top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_right_in[54], chanx_right_in[110], chanx_right_in[166], chanx_left_in[2], chanx_left_in[11], chanx_left_in[58], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size14_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_34_sram_inv[0:7]),
		.out(chany_top_out[160]));

	mux_2level_tapbuf_size14 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_17_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_25_, top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_33_, top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_right_in[0], chanx_right_in[3], chanx_right_in[56], chanx_right_in[112], chanx_left_in[1], chanx_left_in[7], chanx_left_in[57], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size14_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_35_sram_inv[0:7]),
		.out(chany_top_out[164]));

	mux_2level_tapbuf_size14 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[56], chany_top_in[112], chany_bottom_in[54], chany_bottom_in[110], chany_bottom_in[166], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size14_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_36_sram_inv[0:7]),
		.out(chanx_left_out[0]));

	mux_2level_tapbuf_size14 mux_left_track_17 (
		.in({chany_top_in[53], chany_top_in[109], chany_top_in[163], chany_top_in[165], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[57], chany_bottom_in[113], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_}),
		.sram(mux_2level_tapbuf_size14_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_37_sram_inv[0:7]),
		.out(chanx_left_out[8]));

	mux_2level_tapbuf_size14 mux_left_track_25 (
		.in({chany_top_in[52], chany_top_in[108], chany_top_in[159], chany_top_in[164], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[58], chany_bottom_in[114], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_}),
		.sram(mux_2level_tapbuf_size14_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_38_sram_inv[0:7]),
		.out(chanx_left_out[12]));

	mux_2level_tapbuf_size14 mux_left_track_33 (
		.in({chany_top_in[50], chany_top_in[106], chany_top_in[155], chany_top_in[162], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[60], chany_bottom_in[116], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.sram(mux_2level_tapbuf_size14_39_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_39_sram_inv[0:7]),
		.out(chanx_left_out[16]));

	mux_2level_tapbuf_size14 mux_left_track_41 (
		.in({chany_top_in[49], chany_top_in[105], chany_top_in[151], chany_top_in[161], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[61], chany_bottom_in[117], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_}),
		.sram(mux_2level_tapbuf_size14_40_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_40_sram_inv[0:7]),
		.out(chanx_left_out[20]));

	mux_2level_tapbuf_size14 mux_left_track_49 (
		.in({chany_top_in[48], chany_top_in[104], chany_top_in[147], chany_top_in[160], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[62], chany_bottom_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_8_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size14_41_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_41_sram_inv[0:7]),
		.out(chanx_left_out[24]));

	mux_2level_tapbuf_size14 mux_left_track_57 (
		.in({chany_top_in[46], chany_top_in[102], chany_top_in[143], chany_top_in[158], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[64], chany_bottom_in[120], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_42_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_42_sram_inv[0:7]),
		.out(chanx_left_out[28]));

	mux_2level_tapbuf_size14 mux_left_track_73 (
		.in({chany_top_in[44], chany_top_in[100], chany_top_in[135], chany_top_in[156], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[66], chany_bottom_in[122], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_}),
		.sram(mux_2level_tapbuf_size14_43_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_43_sram_inv[0:7]),
		.out(chanx_left_out[36]));

	mux_2level_tapbuf_size14 mux_left_track_81 (
		.in({chany_top_in[42], chany_top_in[98], chany_top_in[131], chany_top_in[154], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[68], chany_bottom_in[124], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_}),
		.sram(mux_2level_tapbuf_size14_44_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_44_sram_inv[0:7]),
		.out(chanx_left_out[40]));

	mux_2level_tapbuf_size14 mux_left_track_89 (
		.in({chany_top_in[41], chany_top_in[97], chany_top_in[127], chany_top_in[153], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[69], chany_bottom_in[125], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_}),
		.sram(mux_2level_tapbuf_size14_45_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_45_sram_inv[0:7]),
		.out(chanx_left_out[44]));

	mux_2level_tapbuf_size14 mux_left_track_97 (
		.in({chany_top_in[40], chany_top_in[96], chany_top_in[123], chany_top_in[152], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[70], chany_bottom_in[126], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.sram(mux_2level_tapbuf_size14_46_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_46_sram_inv[0:7]),
		.out(chanx_left_out[48]));

	mux_2level_tapbuf_size14 mux_left_track_105 (
		.in({chany_top_in[38], chany_top_in[94], chany_top_in[119], chany_top_in[150], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[72], chany_bottom_in[128], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_}),
		.sram(mux_2level_tapbuf_size14_47_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_47_sram_inv[0:7]),
		.out(chanx_left_out[52]));

	mux_2level_tapbuf_size14 mux_left_track_113 (
		.in({chany_top_in[37], chany_top_in[93], chany_top_in[115], chany_top_in[149], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[73], chany_bottom_in[129], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_16_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size14_48_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_48_sram_inv[0:7]),
		.out(chanx_left_out[56]));

	mux_2level_tapbuf_size14 mux_left_track_121 (
		.in({chany_top_in[36], chany_top_in[92], chany_top_in[111], chany_top_in[148], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[74], chany_bottom_in[130], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_49_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_49_sram_inv[0:7]),
		.out(chanx_left_out[60]));

	mux_2level_tapbuf_size14 mux_left_track_137 (
		.in({chany_top_in[33], chany_top_in[89], chany_top_in[103], chany_top_in[145], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[77], chany_bottom_in[133], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_}),
		.sram(mux_2level_tapbuf_size14_50_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_50_sram_inv[0:7]),
		.out(chanx_left_out[68]));

	mux_2level_tapbuf_size14 mux_left_track_145 (
		.in({chany_top_in[32], chany_top_in[88], chany_top_in[99], chany_top_in[144], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[78], chany_bottom_in[134], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_}),
		.sram(mux_2level_tapbuf_size14_51_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_51_sram_inv[0:7]),
		.out(chanx_left_out[72]));

	mux_2level_tapbuf_size14 mux_left_track_153 (
		.in({chany_top_in[30], chany_top_in[86], chany_top_in[95], chany_top_in[142], chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[80], chany_bottom_in[136], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_}),
		.sram(mux_2level_tapbuf_size14_52_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_52_sram_inv[0:7]),
		.out(chanx_left_out[76]));

	mux_2level_tapbuf_size14 mux_left_track_161 (
		.in({chany_top_in[29], chany_top_in[85], chany_top_in[91], chany_top_in[141], chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[81], chany_bottom_in[137], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.sram(mux_2level_tapbuf_size14_53_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_53_sram_inv[0:7]),
		.out(chanx_left_out[80]));

	mux_2level_tapbuf_size14 mux_left_track_169 (
		.in({chany_top_in[28], chany_top_in[84], chany_top_in[87], chany_top_in[140], chany_bottom_in[26], chany_bottom_in[82:83], chany_bottom_in[138], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_}),
		.sram(mux_2level_tapbuf_size14_54_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_54_sram_inv[0:7]),
		.out(chanx_left_out[84]));

	mux_2level_tapbuf_size14 mux_left_track_177 (
		.in({chany_top_in[26], chany_top_in[82:83], chany_top_in[138], chany_bottom_in[28], chany_bottom_in[84], chany_bottom_in[87], chany_bottom_in[140], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_24_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size14_55_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_55_sram_inv[0:7]),
		.out(chanx_left_out[88]));

	mux_2level_tapbuf_size14 mux_left_track_185 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[81], chany_top_in[137], chany_bottom_in[29], chany_bottom_in[85], chany_bottom_in[91], chany_bottom_in[141], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_56_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_56_sram_inv[0:7]),
		.out(chanx_left_out[92]));

	mux_2level_tapbuf_size14 mux_left_track_201 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[78], chany_top_in[134], chany_bottom_in[32], chany_bottom_in[88], chany_bottom_in[99], chany_bottom_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_}),
		.sram(mux_2level_tapbuf_size14_57_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_57_sram_inv[0:7]),
		.out(chanx_left_out[100]));

	mux_2level_tapbuf_size14 mux_left_track_209 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[77], chany_top_in[133], chany_bottom_in[33], chany_bottom_in[89], chany_bottom_in[103], chany_bottom_in[145], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_}),
		.sram(mux_2level_tapbuf_size14_58_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_58_sram_inv[0:7]),
		.out(chanx_left_out[104]));

	mux_2level_tapbuf_size14 mux_left_track_217 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[76], chany_top_in[132], chany_bottom_in[34], chany_bottom_in[90], chany_bottom_in[107], chany_bottom_in[146], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_}),
		.sram(mux_2level_tapbuf_size14_59_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_59_sram_inv[0:7]),
		.out(chanx_left_out[108]));

	mux_2level_tapbuf_size14 mux_left_track_225 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[74], chany_top_in[130], chany_bottom_in[36], chany_bottom_in[92], chany_bottom_in[111], chany_bottom_in[148], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.sram(mux_2level_tapbuf_size14_60_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_60_sram_inv[0:7]),
		.out(chanx_left_out[112]));

	mux_2level_tapbuf_size14 mux_left_track_233 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[73], chany_top_in[129], chany_bottom_in[37], chany_bottom_in[93], chany_bottom_in[115], chany_bottom_in[149], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_}),
		.sram(mux_2level_tapbuf_size14_61_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_61_sram_inv[0:7]),
		.out(chanx_left_out[116]));

	mux_2level_tapbuf_size14 mux_left_track_241 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[72], chany_top_in[128], chany_bottom_in[38], chany_bottom_in[94], chany_bottom_in[119], chany_bottom_in[150], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_32_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size14_62_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_62_sram_inv[0:7]),
		.out(chanx_left_out[120]));

	mux_2level_tapbuf_size14 mux_left_track_249 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[70], chany_top_in[126], chany_bottom_in[40], chany_bottom_in[96], chany_bottom_in[123], chany_bottom_in[152], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_63_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_63_sram_inv[0:7]),
		.out(chanx_left_out[124]));

	mux_2level_tapbuf_size14 mux_left_track_265 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[68], chany_top_in[124], chany_bottom_in[42], chany_bottom_in[98], chany_bottom_in[131], chany_bottom_in[154], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_}),
		.sram(mux_2level_tapbuf_size14_64_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_64_sram_inv[0:7]),
		.out(chanx_left_out[132]));

	mux_2level_tapbuf_size14 mux_left_track_273 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[66], chany_top_in[122], chany_bottom_in[44], chany_bottom_in[100], chany_bottom_in[135], chany_bottom_in[156], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_}),
		.sram(mux_2level_tapbuf_size14_65_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_65_sram_inv[0:7]),
		.out(chanx_left_out[136]));

	mux_2level_tapbuf_size14 mux_left_track_281 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[65], chany_top_in[121], chany_bottom_in[45], chany_bottom_in[101], chany_bottom_in[139], chany_bottom_in[157], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_3_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_11_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_19_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_27_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_}),
		.sram(mux_2level_tapbuf_size14_66_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_66_sram_inv[0:7]),
		.out(chanx_left_out[140]));

	mux_2level_tapbuf_size14 mux_left_track_289 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[64], chany_top_in[120], chany_bottom_in[46], chany_bottom_in[102], chany_bottom_in[143], chany_bottom_in[158], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_4_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_12_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_20_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_28_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.sram(mux_2level_tapbuf_size14_67_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_67_sram_inv[0:7]),
		.out(chanx_left_out[144]));

	mux_2level_tapbuf_size14 mux_left_track_297 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[62], chany_top_in[118], chany_bottom_in[48], chany_bottom_in[104], chany_bottom_in[147], chany_bottom_in[160], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_5_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_13_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_21_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_29_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_}),
		.sram(mux_2level_tapbuf_size14_68_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_68_sram_inv[0:7]),
		.out(chanx_left_out[148]));

	mux_2level_tapbuf_size14 mux_left_track_305 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[61], chany_top_in[117], chany_bottom_in[49], chany_bottom_in[105], chany_bottom_in[151], chany_bottom_in[161], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size14_69_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_69_sram_inv[0:7]),
		.out(chanx_left_out[152]));

	mux_2level_tapbuf_size14 mux_left_track_313 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[60], chany_top_in[116], chany_bottom_in[50], chany_bottom_in[106], chany_bottom_in[155], chany_bottom_in[162], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_7_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_15_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_23_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_31_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_0_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_70_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_70_sram_inv[0:7]),
		.out(chanx_left_out[156]));

	mux_2level_tapbuf_size14 mux_left_track_329 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[57], chany_top_in[113], chany_bottom_in[53], chany_bottom_in[109], chany_bottom_in[163], chany_bottom_in[165], left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_1_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_9_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_17_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_25_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_33_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size14_71_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size14_71_sram_inv[0:7]),
		.out(chanx_left_out[164]));

	mux_2level_tapbuf_size14_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_0_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_1_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_2_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_3_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_4_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_5_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_6_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_7_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_8_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_9_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_10_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_11_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_12_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_13_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_14_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_15_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_16_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_17_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_18_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_19_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_20_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_21_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_22_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_23_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_24_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_25_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_26_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_27_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_28_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_29_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_30_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_31_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_32_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_33_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_34_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_top_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_35_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_36_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_37_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_38_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_39_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_39_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_40_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_40_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_41_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_41_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_42_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_42_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_43_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_43_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_44_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_44_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_45_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_45_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_46_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_46_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_47_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_47_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_48_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_48_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_49_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_49_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_50_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_50_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_51_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_51_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_52_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_52_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_53_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_53_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_54_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_54_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_55_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_55_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_56_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_56_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_57_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_57_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_58_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_58_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_59_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_59_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_60_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_60_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_61_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_61_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_62_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_62_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_63_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_63_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_64_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_64_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_65_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_65_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_66_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_66_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_67_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_67_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_68_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_68_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_305 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_69_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_69_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_313 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size14_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_70_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_70_sram_inv[0:7]));

	mux_2level_tapbuf_size14_mem mem_left_track_329 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_9_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size14_71_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size14_71_sram_inv[0:7]));

	mux_2level_tapbuf_size7 mux_right_track_0 (
		.in({chany_top_in[54], chany_top_in[110], chany_top_in[166], chany_bottom_in[53], chany_bottom_in[109], chany_bottom_in[163], chany_bottom_in[165]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size7 mux_right_track_328 (
		.in({chany_top_in[53], chany_top_in[109], chany_top_in[163], chany_top_in[165], chany_bottom_in[54], chany_bottom_in[110], chany_bottom_in[166]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chanx_right_out[164]));

	mux_2level_tapbuf_size7 mux_bottom_track_321 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[56], chanx_right_in[112], chanx_left_in[54], chanx_left_in[110], chanx_left_in[166]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chany_bottom_out[160]));

	mux_2level_tapbuf_size7 mux_bottom_track_329 (
		.in({chanx_right_in[54], chanx_right_in[110], chanx_right_in[166], chanx_left_in[0], chanx_left_in[3], chanx_left_in[56], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chany_bottom_out[164]));

	mux_2level_tapbuf_size7_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size14_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_right_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_321 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_329 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[56], chany_top_in[112], chany_bottom_in[52], chany_bottom_in[108], chany_bottom_in[159], chany_bottom_in[164]}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size8 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[57], chany_top_in[113], chany_bottom_in[50], chany_bottom_in[106], chany_bottom_in[155], chany_bottom_in[162]}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size8 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[58], chany_top_in[114], chany_bottom_in[49], chany_bottom_in[105], chany_bottom_in[151], chany_bottom_in[161]}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size8 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[60], chany_top_in[116], chany_bottom_in[48], chany_bottom_in[104], chany_bottom_in[147], chany_bottom_in[160]}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size8 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[61], chany_top_in[117], chany_bottom_in[46], chany_bottom_in[102], chany_bottom_in[143], chany_bottom_in[158]}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size8 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[62], chany_top_in[118], chany_bottom_in[45], chany_bottom_in[101], chany_bottom_in[139], chany_bottom_in[157]}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size8 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[64], chany_top_in[120], chany_bottom_in[44], chany_bottom_in[100], chany_bottom_in[135], chany_bottom_in[156]}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size8 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[65], chany_top_in[121], chany_bottom_in[42], chany_bottom_in[98], chany_bottom_in[131], chany_bottom_in[154]}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size8 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[66], chany_top_in[122], chany_bottom_in[41], chany_bottom_in[97], chany_bottom_in[127], chany_bottom_in[153]}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size8 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[68], chany_top_in[124], chany_bottom_in[40], chany_bottom_in[96], chany_bottom_in[123], chany_bottom_in[152]}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size8 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[69], chany_top_in[125], chany_bottom_in[38], chany_bottom_in[94], chany_bottom_in[119], chany_bottom_in[150]}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size8 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[70], chany_top_in[126], chany_bottom_in[37], chany_bottom_in[93], chany_bottom_in[115], chany_bottom_in[149]}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size8 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[72], chany_top_in[128], chany_bottom_in[36], chany_bottom_in[92], chany_bottom_in[111], chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size8 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[73], chany_top_in[129], chany_bottom_in[34], chany_bottom_in[90], chany_bottom_in[107], chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size8 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[74], chany_top_in[130], chany_bottom_in[33], chany_bottom_in[89], chany_bottom_in[103], chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size8 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[76], chany_top_in[132], chany_bottom_in[32], chany_bottom_in[88], chany_bottom_in[99], chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size8 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[77], chany_top_in[133], chany_bottom_in[30], chany_bottom_in[86], chany_bottom_in[95], chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size8_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_16_sram_inv[0:5]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size8 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[78], chany_top_in[134], chany_bottom_in[29], chany_bottom_in[85], chany_bottom_in[91], chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size8_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_17_sram_inv[0:5]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size8 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[80], chany_top_in[136], chany_bottom_in[28], chany_bottom_in[84], chany_bottom_in[87], chany_bottom_in[140]}),
		.sram(mux_2level_tapbuf_size8_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_18_sram_inv[0:5]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size8 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[81], chany_top_in[137], chany_bottom_in[26], chany_bottom_in[82:83], chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size8_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_19_sram_inv[0:5]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size8 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[82:83], chany_top_in[138], chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[81], chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size8_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_20_sram_inv[0:5]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size8 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[84], chany_top_in[87], chany_top_in[140], chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[80], chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size8_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_21_sram_inv[0:5]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size8 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[85], chany_top_in[91], chany_top_in[141], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[78], chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size8_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_22_sram_inv[0:5]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size8 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[86], chany_top_in[95], chany_top_in[142], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[77], chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size8_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_23_sram_inv[0:5]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size8 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[88], chany_top_in[99], chany_top_in[144], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[76], chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size8_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_24_sram_inv[0:5]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size8 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[89], chany_top_in[103], chany_top_in[145], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[74], chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size8_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_25_sram_inv[0:5]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size8 mux_right_track_216 (
		.in({chany_top_in[34], chany_top_in[90], chany_top_in[107], chany_top_in[146], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[73], chany_bottom_in[129]}),
		.sram(mux_2level_tapbuf_size8_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_26_sram_inv[0:5]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size8 mux_right_track_224 (
		.in({chany_top_in[36], chany_top_in[92], chany_top_in[111], chany_top_in[148], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[72], chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size8_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_27_sram_inv[0:5]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size8 mux_right_track_232 (
		.in({chany_top_in[37], chany_top_in[93], chany_top_in[115], chany_top_in[149], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[70], chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size8_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_28_sram_inv[0:5]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size8 mux_right_track_240 (
		.in({chany_top_in[38], chany_top_in[94], chany_top_in[119], chany_top_in[150], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[69], chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size8_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_29_sram_inv[0:5]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size8 mux_right_track_248 (
		.in({chany_top_in[40], chany_top_in[96], chany_top_in[123], chany_top_in[152], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[68], chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size8_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_30_sram_inv[0:5]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size8 mux_right_track_256 (
		.in({chany_top_in[41], chany_top_in[97], chany_top_in[127], chany_top_in[153], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[66], chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size8_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_31_sram_inv[0:5]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size8 mux_right_track_264 (
		.in({chany_top_in[42], chany_top_in[98], chany_top_in[131], chany_top_in[154], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[65], chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size8_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_32_sram_inv[0:5]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size8 mux_right_track_272 (
		.in({chany_top_in[44], chany_top_in[100], chany_top_in[135], chany_top_in[156], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[64], chany_bottom_in[120]}),
		.sram(mux_2level_tapbuf_size8_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_33_sram_inv[0:5]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size8 mux_right_track_280 (
		.in({chany_top_in[45], chany_top_in[101], chany_top_in[139], chany_top_in[157], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[62], chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size8_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_34_sram_inv[0:5]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size8 mux_right_track_288 (
		.in({chany_top_in[46], chany_top_in[102], chany_top_in[143], chany_top_in[158], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[61], chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size8_35_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_35_sram_inv[0:5]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size8 mux_right_track_296 (
		.in({chany_top_in[48], chany_top_in[104], chany_top_in[147], chany_top_in[160], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[60], chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size8_36_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_36_sram_inv[0:5]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size8 mux_right_track_304 (
		.in({chany_top_in[49], chany_top_in[105], chany_top_in[151], chany_top_in[161], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[58], chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size8_37_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_37_sram_inv[0:5]),
		.out(chanx_right_out[152]));

	mux_2level_tapbuf_size8 mux_right_track_312 (
		.in({chany_top_in[50], chany_top_in[106], chany_top_in[155], chany_top_in[162], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[57], chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size8_38_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_38_sram_inv[0:5]),
		.out(chanx_right_out[156]));

	mux_2level_tapbuf_size8 mux_right_track_320 (
		.in({chany_top_in[52], chany_top_in[108], chany_top_in[159], chany_top_in[164], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[56], chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size8_39_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_39_sram_inv[0:5]),
		.out(chanx_right_out[160]));

	mux_2level_tapbuf_size8 mux_bottom_track_1 (
		.in({chanx_right_in[53], chanx_right_in[109], chanx_right_in[163], chanx_right_in[165], chanx_left_in[1], chanx_left_in[7], chanx_left_in[57], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size8_40_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_40_sram_inv[0:5]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size8 mux_bottom_track_9 (
		.in({chanx_right_in[52], chanx_right_in[108], chanx_right_in[159], chanx_right_in[164], chanx_left_in[2], chanx_left_in[11], chanx_left_in[58], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size8_41_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_41_sram_inv[0:5]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size8 mux_bottom_track_17 (
		.in({chanx_right_in[50], chanx_right_in[106], chanx_right_in[155], chanx_right_in[162], chanx_left_in[4], chanx_left_in[15], chanx_left_in[60], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size8_42_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_42_sram_inv[0:5]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size8 mux_bottom_track_25 (
		.in({chanx_right_in[49], chanx_right_in[105], chanx_right_in[151], chanx_right_in[161], chanx_left_in[5], chanx_left_in[19], chanx_left_in[61], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size8_43_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_43_sram_inv[0:5]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size8 mux_bottom_track_33 (
		.in({chanx_right_in[48], chanx_right_in[104], chanx_right_in[147], chanx_right_in[160], chanx_left_in[6], chanx_left_in[23], chanx_left_in[62], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size8_44_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_44_sram_inv[0:5]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size8 mux_bottom_track_41 (
		.in({chanx_right_in[46], chanx_right_in[102], chanx_right_in[143], chanx_right_in[158], chanx_left_in[8], chanx_left_in[27], chanx_left_in[64], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size8_45_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_45_sram_inv[0:5]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size8 mux_bottom_track_49 (
		.in({chanx_right_in[45], chanx_right_in[101], chanx_right_in[139], chanx_right_in[157], chanx_left_in[9], chanx_left_in[31], chanx_left_in[65], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size8_46_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_46_sram_inv[0:5]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size8 mux_bottom_track_57 (
		.in({chanx_right_in[44], chanx_right_in[100], chanx_right_in[135], chanx_right_in[156], chanx_left_in[10], chanx_left_in[35], chanx_left_in[66], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size8_47_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_47_sram_inv[0:5]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size8 mux_bottom_track_65 (
		.in({chanx_right_in[42], chanx_right_in[98], chanx_right_in[131], chanx_right_in[154], chanx_left_in[12], chanx_left_in[39], chanx_left_in[68], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size8_48_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_48_sram_inv[0:5]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size8 mux_bottom_track_73 (
		.in({chanx_right_in[41], chanx_right_in[97], chanx_right_in[127], chanx_right_in[153], chanx_left_in[13], chanx_left_in[43], chanx_left_in[69], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size8_49_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_49_sram_inv[0:5]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size8 mux_bottom_track_81 (
		.in({chanx_right_in[40], chanx_right_in[96], chanx_right_in[123], chanx_right_in[152], chanx_left_in[14], chanx_left_in[47], chanx_left_in[70], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size8_50_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_50_sram_inv[0:5]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size8 mux_bottom_track_89 (
		.in({chanx_right_in[38], chanx_right_in[94], chanx_right_in[119], chanx_right_in[150], chanx_left_in[16], chanx_left_in[51], chanx_left_in[72], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size8_51_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_51_sram_inv[0:5]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size8 mux_bottom_track_97 (
		.in({chanx_right_in[37], chanx_right_in[93], chanx_right_in[115], chanx_right_in[149], chanx_left_in[17], chanx_left_in[55], chanx_left_in[73], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size8_52_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_52_sram_inv[0:5]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size8 mux_bottom_track_105 (
		.in({chanx_right_in[36], chanx_right_in[92], chanx_right_in[111], chanx_right_in[148], chanx_left_in[18], chanx_left_in[59], chanx_left_in[74], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size8_53_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_53_sram_inv[0:5]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size8 mux_bottom_track_113 (
		.in({chanx_right_in[34], chanx_right_in[90], chanx_right_in[107], chanx_right_in[146], chanx_left_in[20], chanx_left_in[63], chanx_left_in[76], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size8_54_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_54_sram_inv[0:5]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size8 mux_bottom_track_121 (
		.in({chanx_right_in[33], chanx_right_in[89], chanx_right_in[103], chanx_right_in[145], chanx_left_in[21], chanx_left_in[67], chanx_left_in[77], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size8_55_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_55_sram_inv[0:5]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size8 mux_bottom_track_129 (
		.in({chanx_right_in[32], chanx_right_in[88], chanx_right_in[99], chanx_right_in[144], chanx_left_in[22], chanx_left_in[71], chanx_left_in[78], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size8_56_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_56_sram_inv[0:5]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size8 mux_bottom_track_137 (
		.in({chanx_right_in[30], chanx_right_in[86], chanx_right_in[95], chanx_right_in[142], chanx_left_in[24], chanx_left_in[75], chanx_left_in[80], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size8_57_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_57_sram_inv[0:5]),
		.out(chany_bottom_out[68]));

	mux_2level_tapbuf_size8 mux_bottom_track_145 (
		.in({chanx_right_in[29], chanx_right_in[85], chanx_right_in[91], chanx_right_in[141], chanx_left_in[25], chanx_left_in[79], chanx_left_in[81], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size8_58_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_58_sram_inv[0:5]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size8 mux_bottom_track_153 (
		.in({chanx_right_in[28], chanx_right_in[84], chanx_right_in[87], chanx_right_in[140], chanx_left_in[26], chanx_left_in[82:83], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size8_59_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_59_sram_inv[0:5]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size8 mux_bottom_track_161 (
		.in({chanx_right_in[26], chanx_right_in[82:83], chanx_right_in[138], chanx_left_in[28], chanx_left_in[84], chanx_left_in[87], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size8_60_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_60_sram_inv[0:5]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size8 mux_bottom_track_169 (
		.in({chanx_right_in[25], chanx_right_in[79], chanx_right_in[81], chanx_right_in[137], chanx_left_in[29], chanx_left_in[85], chanx_left_in[91], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size8_61_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_61_sram_inv[0:5]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size8 mux_bottom_track_177 (
		.in({chanx_right_in[24], chanx_right_in[75], chanx_right_in[80], chanx_right_in[136], chanx_left_in[30], chanx_left_in[86], chanx_left_in[95], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size8_62_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_62_sram_inv[0:5]),
		.out(chany_bottom_out[88]));

	mux_2level_tapbuf_size8 mux_bottom_track_185 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[78], chanx_right_in[134], chanx_left_in[32], chanx_left_in[88], chanx_left_in[99], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size8_63_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_63_sram_inv[0:5]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size8 mux_bottom_track_193 (
		.in({chanx_right_in[21], chanx_right_in[67], chanx_right_in[77], chanx_right_in[133], chanx_left_in[33], chanx_left_in[89], chanx_left_in[103], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size8_64_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_64_sram_inv[0:5]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size8 mux_bottom_track_201 (
		.in({chanx_right_in[20], chanx_right_in[63], chanx_right_in[76], chanx_right_in[132], chanx_left_in[34], chanx_left_in[90], chanx_left_in[107], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size8_65_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_65_sram_inv[0:5]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size8 mux_bottom_track_209 (
		.in({chanx_right_in[18], chanx_right_in[59], chanx_right_in[74], chanx_right_in[130], chanx_left_in[36], chanx_left_in[92], chanx_left_in[111], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size8_66_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_66_sram_inv[0:5]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size8 mux_bottom_track_217 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[73], chanx_right_in[129], chanx_left_in[37], chanx_left_in[93], chanx_left_in[115], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size8_67_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_67_sram_inv[0:5]),
		.out(chany_bottom_out[108]));

	mux_2level_tapbuf_size8 mux_bottom_track_225 (
		.in({chanx_right_in[16], chanx_right_in[51], chanx_right_in[72], chanx_right_in[128], chanx_left_in[38], chanx_left_in[94], chanx_left_in[119], chanx_left_in[150]}),
		.sram(mux_2level_tapbuf_size8_68_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_68_sram_inv[0:5]),
		.out(chany_bottom_out[112]));

	mux_2level_tapbuf_size8 mux_bottom_track_233 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[70], chanx_right_in[126], chanx_left_in[40], chanx_left_in[96], chanx_left_in[123], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size8_69_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_69_sram_inv[0:5]),
		.out(chany_bottom_out[116]));

	mux_2level_tapbuf_size8 mux_bottom_track_241 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[69], chanx_right_in[125], chanx_left_in[41], chanx_left_in[97], chanx_left_in[127], chanx_left_in[153]}),
		.sram(mux_2level_tapbuf_size8_70_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_70_sram_inv[0:5]),
		.out(chany_bottom_out[120]));

	mux_2level_tapbuf_size8 mux_bottom_track_249 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[68], chanx_right_in[124], chanx_left_in[42], chanx_left_in[98], chanx_left_in[131], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size8_71_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_71_sram_inv[0:5]),
		.out(chany_bottom_out[124]));

	mux_2level_tapbuf_size8 mux_bottom_track_257 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[66], chanx_right_in[122], chanx_left_in[44], chanx_left_in[100], chanx_left_in[135], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size8_72_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_72_sram_inv[0:5]),
		.out(chany_bottom_out[128]));

	mux_2level_tapbuf_size8 mux_bottom_track_265 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[65], chanx_right_in[121], chanx_left_in[45], chanx_left_in[101], chanx_left_in[139], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size8_73_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_73_sram_inv[0:5]),
		.out(chany_bottom_out[132]));

	mux_2level_tapbuf_size8 mux_bottom_track_273 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[64], chanx_right_in[120], chanx_left_in[46], chanx_left_in[102], chanx_left_in[143], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size8_74_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_74_sram_inv[0:5]),
		.out(chany_bottom_out[136]));

	mux_2level_tapbuf_size8 mux_bottom_track_281 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[62], chanx_right_in[118], chanx_left_in[48], chanx_left_in[104], chanx_left_in[147], chanx_left_in[160]}),
		.sram(mux_2level_tapbuf_size8_75_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_75_sram_inv[0:5]),
		.out(chany_bottom_out[140]));

	mux_2level_tapbuf_size8 mux_bottom_track_289 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[61], chanx_right_in[117], chanx_left_in[49], chanx_left_in[105], chanx_left_in[151], chanx_left_in[161]}),
		.sram(mux_2level_tapbuf_size8_76_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_76_sram_inv[0:5]),
		.out(chany_bottom_out[144]));

	mux_2level_tapbuf_size8 mux_bottom_track_297 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[60], chanx_right_in[116], chanx_left_in[50], chanx_left_in[106], chanx_left_in[155], chanx_left_in[162]}),
		.sram(mux_2level_tapbuf_size8_77_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_77_sram_inv[0:5]),
		.out(chany_bottom_out[148]));

	mux_2level_tapbuf_size8 mux_bottom_track_305 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[58], chanx_right_in[114], chanx_left_in[52], chanx_left_in[108], chanx_left_in[159], chanx_left_in[164]}),
		.sram(mux_2level_tapbuf_size8_78_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_78_sram_inv[0:5]),
		.out(chany_bottom_out[152]));

	mux_2level_tapbuf_size8 mux_bottom_track_313 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[57], chanx_right_in[113], chanx_left_in[53], chanx_left_in[109], chanx_left_in[163], chanx_left_in[165]}),
		.sram(mux_2level_tapbuf_size8_79_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_79_sram_inv[0:5]),
		.out(chany_bottom_out[156]));

	mux_2level_tapbuf_size8_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_16_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_17_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_18_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_19_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_20_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_21_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_22_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_23_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_24_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_25_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_26_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_27_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_28_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_29_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_30_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_31_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_32_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_33_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_34_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_35_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_35_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_36_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_36_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_37_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_37_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_38_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_38_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_right_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_39_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_39_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_40_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_40_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_41_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_41_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_42_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_42_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_43_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_43_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_44_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_44_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_45_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_45_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_46_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_46_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_47_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_47_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_48_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_48_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_49_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_49_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_50_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_50_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_51_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_51_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_52_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_52_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_53_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_53_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_54_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_54_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_55_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_55_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_56_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_56_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_57_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_57_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_58_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_58_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_59_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_59_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_60_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_60_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_61_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_61_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_62_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_62_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_63_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_63_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_64_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_64_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_65_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_65_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_66_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_66_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_67_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_67_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_68_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_68_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_69_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_69_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_70_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_70_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_71_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_71_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_72_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_72_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_73_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_73_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_74_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_74_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_75_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_75_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_76_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_76_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_77_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_77_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_305 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_78_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_78_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_313 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_79_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_79_sram_inv[0:5]));

endmodule
// ----- END Verilog module for sb_3__2_ -----

//----- Default net type -----
`default_nettype wire



