module router_bench (
    input   [34:0] idata_0,
    input              ivalid_0, 
    input      ivch_0,   
    output   [1:0]   oack_0 ,   
    output   [1:0]   ordy_0 ,   
    output   [1:0]   olck_0 ,   
    input   [34:0] idata_1 ,
    input              ivalid_1 ,
    input      ivch_1 ,
    output   [1:0]   oack_1 ,
    output   [1:0]   ordy_1 ,
    output   [1:0]   olck_1 ,
    input   [34:0] idata_2 ,
    input              ivalid_2 , 
    input      ivch_2 ,
    output   [1:0]   oack_2 ,  
    output   [1:0]   ordy_2 ,  
    output   [1:0]   olck_2 ,  
    input   [34:0] idata_3 ,  
    input              ivalid_3 , 
    input      ivch_3 ,   
    output   [1:0]   oack_3 ,   
    output   [1:0]   ordy_3 ,   
    output   [1:0]   olck_3 ,   
    input   [34:0] idata_4 ,  
    input              ivalid_4 , 
    input      ivch_4 ,   
    output   [1:0]   oack_4 ,   
    output   [1:0]   ordy_4 ,   
    output   [1:0]   olck_4 ,   
    output   [34:0] odata_0 , 
    output            ovalid_0 ,
    output      ovch_0 ,   
    input   [1:0]   iack_0 , 
    input   [1:0]   ilck_0 ,
    output   [34:0] odata_1 ,
    output              ovalid_1 , 
    output      ovch_1 ,
    input   [1:0]   iack_1 ,   
    input   [1:0]   ilck_1 ,   
    output   [34:0] odata_2 ,
    output              ovalid_2 ,
    output      ovch_2 ,
    input   [1:0]   iack_2 ,
    input   [1:0]   ilck_2 ,
    output   [34:0] odata_3 ,
    output              ovalid_3 , 
    output      ovch_3 ,   
    input   [1:0]   iack_3 ,   
    input   [1:0]   ilck_3 ,   
    output   [34:0] odata_4 , 
    output              ovalid_4 , 
    output      ovch_4 ,   
    input   [1:0]   iack_4 ,   
    input   [1:0]   ilck_4 ,   
    input [1:0]  my_xpos ,
    input [1:0]  my_ypos ,

    input    clk ,
    input    rst_    );

router rtr0 ( 

    .oack_0(oack_0) ,
    .ordy_0(ordy_0) ,
    .olck_0(olck_0) ,
    .oack_1(oack_1) ,
    .ordy_1(ordy_1) ,
    .olck_1(olck_1) ,
    .oack_2(oack_2) ,
    .ordy_2(ordy_2) ,
    .olck_2(olck_2) ,
    .oack_3(oack_3) ,
    .ordy_3(ordy_3) ,
    .olck_3(olck_3) ,
    .oack_4(oack_4) ,
    .ordy_4(ordy_4) ,
    .olck_4(olck_4) ,
    .odata_0(odata_0) ,
    .ovalid_0(ovalid_0) ,
    .ovch_0(ovch_0) ,
    .odata_1(odata_1) ,
    .ovalid_1(ovalid_1) ,
    .ovch_1(ovch_1) ,
    .odata_2(odata_2) ,
    .ovalid_2(ovalid_2) ,
    .ovch_2(ovch_2) ,
    .odata_3(odata_3) ,
    .ovalid_3(ovalid_3) ,
    .ovch_3(ovch_3) ,
    .odata_4(odata_4) ,
    .ovalid_4(ovalid_4) ,
    .ovch_4(ovch_4) ,
    .idata_0(idata_0) ,
    .ivalid_0(ivalid_0) ,
    .ivch_0(ivch_0) ,
    .idata_1(idata_1) ,
    .ivalid_1(ivalid_1) ,
    .ivch_1(ivch_1) ,
    .idata_2(idata_2) ,
    .ivalid_2(ivalid_2) ,
    .ivch_2(ivch_2) ,
    .idata_3(idata_3) ,
    .ivalid_3(ivalid_3) ,
    .ivch_3(ivch_3) ,
    .idata_4(idata_4) ,
    .ivalid_4(ivalid_4) ,
    .ivch_4(ivch_4) ,
    .iack_0(iack_0) ,
    .ilck_0(ilck_0) ,
    .iack_1(iack_1) ,
    .ilck_1(ilck_1) ,
    .iack_2(iack_2) ,
    .ilck_2(ilck_2) ,
    .iack_3(iack_3) ,
    .ilck_3(ilck_3) ,
    .iack_4(iack_4) ,
    .ilck_4(ilck_4) ,
    .my_xpos(my_xpos) ,
    .my_ypos(my_ypos) ,
    .clk(clk) ,
    .rst_(rst_) 

); 

endmodule

       

