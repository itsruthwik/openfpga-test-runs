//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Oct 17 11:38:19 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__2_ -----
module sb_0__2_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:159] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:159] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:159] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:159] chany_top_out;
//----- OUTPUT PORTS -----
output [0:159] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:159] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size10_0_sram;
wire [0:7] mux_2level_tapbuf_size10_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_10_sram;
wire [0:7] mux_2level_tapbuf_size10_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_11_sram;
wire [0:7] mux_2level_tapbuf_size10_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_12_sram;
wire [0:7] mux_2level_tapbuf_size10_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_13_sram;
wire [0:7] mux_2level_tapbuf_size10_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_14_sram;
wire [0:7] mux_2level_tapbuf_size10_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_15_sram;
wire [0:7] mux_2level_tapbuf_size10_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_16_sram;
wire [0:7] mux_2level_tapbuf_size10_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_17_sram;
wire [0:7] mux_2level_tapbuf_size10_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_18_sram;
wire [0:7] mux_2level_tapbuf_size10_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_19_sram;
wire [0:7] mux_2level_tapbuf_size10_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_1_sram;
wire [0:7] mux_2level_tapbuf_size10_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_20_sram;
wire [0:7] mux_2level_tapbuf_size10_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_21_sram;
wire [0:7] mux_2level_tapbuf_size10_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_22_sram;
wire [0:7] mux_2level_tapbuf_size10_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_23_sram;
wire [0:7] mux_2level_tapbuf_size10_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_24_sram;
wire [0:7] mux_2level_tapbuf_size10_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_25_sram;
wire [0:7] mux_2level_tapbuf_size10_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_26_sram;
wire [0:7] mux_2level_tapbuf_size10_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_27_sram;
wire [0:7] mux_2level_tapbuf_size10_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_28_sram;
wire [0:7] mux_2level_tapbuf_size10_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_29_sram;
wire [0:7] mux_2level_tapbuf_size10_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_2_sram;
wire [0:7] mux_2level_tapbuf_size10_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_30_sram;
wire [0:7] mux_2level_tapbuf_size10_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_31_sram;
wire [0:7] mux_2level_tapbuf_size10_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_3_sram;
wire [0:7] mux_2level_tapbuf_size10_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_4_sram;
wire [0:7] mux_2level_tapbuf_size10_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_5_sram;
wire [0:7] mux_2level_tapbuf_size10_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_6_sram;
wire [0:7] mux_2level_tapbuf_size10_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_7_sram;
wire [0:7] mux_2level_tapbuf_size10_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_8_sram;
wire [0:7] mux_2level_tapbuf_size10_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size10_9_sram;
wire [0:7] mux_2level_tapbuf_size10_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size10_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size11_0_sram;
wire [0:7] mux_2level_tapbuf_size11_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_1_sram;
wire [0:7] mux_2level_tapbuf_size11_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_2_sram;
wire [0:7] mux_2level_tapbuf_size11_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_3_sram;
wire [0:7] mux_2level_tapbuf_size11_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_4_sram;
wire [0:7] mux_2level_tapbuf_size11_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_5_sram;
wire [0:7] mux_2level_tapbuf_size11_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_6_sram;
wire [0:7] mux_2level_tapbuf_size11_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_7_sram;
wire [0:7] mux_2level_tapbuf_size11_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_8_sram;
wire [0:7] mux_2level_tapbuf_size11_8_sram_inv;
wire [0:0] mux_2level_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_8_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_100_sram;
wire [0:1] mux_2level_tapbuf_size3_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_101_sram;
wire [0:1] mux_2level_tapbuf_size3_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_102_sram;
wire [0:1] mux_2level_tapbuf_size3_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_103_sram;
wire [0:1] mux_2level_tapbuf_size3_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_104_sram;
wire [0:1] mux_2level_tapbuf_size3_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_105_sram;
wire [0:1] mux_2level_tapbuf_size3_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_106_sram;
wire [0:1] mux_2level_tapbuf_size3_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_107_sram;
wire [0:1] mux_2level_tapbuf_size3_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_108_sram;
wire [0:1] mux_2level_tapbuf_size3_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_109_sram;
wire [0:1] mux_2level_tapbuf_size3_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_10_sram;
wire [0:1] mux_2level_tapbuf_size3_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_110_sram;
wire [0:1] mux_2level_tapbuf_size3_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_111_sram;
wire [0:1] mux_2level_tapbuf_size3_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_112_sram;
wire [0:1] mux_2level_tapbuf_size3_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_113_sram;
wire [0:1] mux_2level_tapbuf_size3_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_114_sram;
wire [0:1] mux_2level_tapbuf_size3_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_115_sram;
wire [0:1] mux_2level_tapbuf_size3_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_116_sram;
wire [0:1] mux_2level_tapbuf_size3_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_117_sram;
wire [0:1] mux_2level_tapbuf_size3_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_118_sram;
wire [0:1] mux_2level_tapbuf_size3_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_119_sram;
wire [0:1] mux_2level_tapbuf_size3_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_11_sram;
wire [0:1] mux_2level_tapbuf_size3_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_120_sram;
wire [0:1] mux_2level_tapbuf_size3_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_121_sram;
wire [0:1] mux_2level_tapbuf_size3_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_122_sram;
wire [0:1] mux_2level_tapbuf_size3_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_123_sram;
wire [0:1] mux_2level_tapbuf_size3_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_124_sram;
wire [0:1] mux_2level_tapbuf_size3_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_125_sram;
wire [0:1] mux_2level_tapbuf_size3_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_126_sram;
wire [0:1] mux_2level_tapbuf_size3_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_127_sram;
wire [0:1] mux_2level_tapbuf_size3_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_128_sram;
wire [0:1] mux_2level_tapbuf_size3_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_129_sram;
wire [0:1] mux_2level_tapbuf_size3_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_12_sram;
wire [0:1] mux_2level_tapbuf_size3_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_130_sram;
wire [0:1] mux_2level_tapbuf_size3_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_131_sram;
wire [0:1] mux_2level_tapbuf_size3_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_132_sram;
wire [0:1] mux_2level_tapbuf_size3_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_133_sram;
wire [0:1] mux_2level_tapbuf_size3_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_134_sram;
wire [0:1] mux_2level_tapbuf_size3_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_135_sram;
wire [0:1] mux_2level_tapbuf_size3_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_136_sram;
wire [0:1] mux_2level_tapbuf_size3_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_137_sram;
wire [0:1] mux_2level_tapbuf_size3_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_138_sram;
wire [0:1] mux_2level_tapbuf_size3_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_139_sram;
wire [0:1] mux_2level_tapbuf_size3_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_13_sram;
wire [0:1] mux_2level_tapbuf_size3_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_140_sram;
wire [0:1] mux_2level_tapbuf_size3_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_141_sram;
wire [0:1] mux_2level_tapbuf_size3_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_142_sram;
wire [0:1] mux_2level_tapbuf_size3_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_143_sram;
wire [0:1] mux_2level_tapbuf_size3_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_144_sram;
wire [0:1] mux_2level_tapbuf_size3_144_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_145_sram;
wire [0:1] mux_2level_tapbuf_size3_145_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_146_sram;
wire [0:1] mux_2level_tapbuf_size3_146_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_147_sram;
wire [0:1] mux_2level_tapbuf_size3_147_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_148_sram;
wire [0:1] mux_2level_tapbuf_size3_148_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_149_sram;
wire [0:1] mux_2level_tapbuf_size3_149_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_14_sram;
wire [0:1] mux_2level_tapbuf_size3_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_150_sram;
wire [0:1] mux_2level_tapbuf_size3_150_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_151_sram;
wire [0:1] mux_2level_tapbuf_size3_151_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_152_sram;
wire [0:1] mux_2level_tapbuf_size3_152_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_153_sram;
wire [0:1] mux_2level_tapbuf_size3_153_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_154_sram;
wire [0:1] mux_2level_tapbuf_size3_154_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_155_sram;
wire [0:1] mux_2level_tapbuf_size3_155_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_156_sram;
wire [0:1] mux_2level_tapbuf_size3_156_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_157_sram;
wire [0:1] mux_2level_tapbuf_size3_157_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_158_sram;
wire [0:1] mux_2level_tapbuf_size3_158_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_159_sram;
wire [0:1] mux_2level_tapbuf_size3_159_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_15_sram;
wire [0:1] mux_2level_tapbuf_size3_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_16_sram;
wire [0:1] mux_2level_tapbuf_size3_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_17_sram;
wire [0:1] mux_2level_tapbuf_size3_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_18_sram;
wire [0:1] mux_2level_tapbuf_size3_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_19_sram;
wire [0:1] mux_2level_tapbuf_size3_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_20_sram;
wire [0:1] mux_2level_tapbuf_size3_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_21_sram;
wire [0:1] mux_2level_tapbuf_size3_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_22_sram;
wire [0:1] mux_2level_tapbuf_size3_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_23_sram;
wire [0:1] mux_2level_tapbuf_size3_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_24_sram;
wire [0:1] mux_2level_tapbuf_size3_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_25_sram;
wire [0:1] mux_2level_tapbuf_size3_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_26_sram;
wire [0:1] mux_2level_tapbuf_size3_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_27_sram;
wire [0:1] mux_2level_tapbuf_size3_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_28_sram;
wire [0:1] mux_2level_tapbuf_size3_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_29_sram;
wire [0:1] mux_2level_tapbuf_size3_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_30_sram;
wire [0:1] mux_2level_tapbuf_size3_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_31_sram;
wire [0:1] mux_2level_tapbuf_size3_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_32_sram;
wire [0:1] mux_2level_tapbuf_size3_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_33_sram;
wire [0:1] mux_2level_tapbuf_size3_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_34_sram;
wire [0:1] mux_2level_tapbuf_size3_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_35_sram;
wire [0:1] mux_2level_tapbuf_size3_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_36_sram;
wire [0:1] mux_2level_tapbuf_size3_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_37_sram;
wire [0:1] mux_2level_tapbuf_size3_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_38_sram;
wire [0:1] mux_2level_tapbuf_size3_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_39_sram;
wire [0:1] mux_2level_tapbuf_size3_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_40_sram;
wire [0:1] mux_2level_tapbuf_size3_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_41_sram;
wire [0:1] mux_2level_tapbuf_size3_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_42_sram;
wire [0:1] mux_2level_tapbuf_size3_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_43_sram;
wire [0:1] mux_2level_tapbuf_size3_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_44_sram;
wire [0:1] mux_2level_tapbuf_size3_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_45_sram;
wire [0:1] mux_2level_tapbuf_size3_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_46_sram;
wire [0:1] mux_2level_tapbuf_size3_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_47_sram;
wire [0:1] mux_2level_tapbuf_size3_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_48_sram;
wire [0:1] mux_2level_tapbuf_size3_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_49_sram;
wire [0:1] mux_2level_tapbuf_size3_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_50_sram;
wire [0:1] mux_2level_tapbuf_size3_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_51_sram;
wire [0:1] mux_2level_tapbuf_size3_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_52_sram;
wire [0:1] mux_2level_tapbuf_size3_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_53_sram;
wire [0:1] mux_2level_tapbuf_size3_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_54_sram;
wire [0:1] mux_2level_tapbuf_size3_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_55_sram;
wire [0:1] mux_2level_tapbuf_size3_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_56_sram;
wire [0:1] mux_2level_tapbuf_size3_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_57_sram;
wire [0:1] mux_2level_tapbuf_size3_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_58_sram;
wire [0:1] mux_2level_tapbuf_size3_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_59_sram;
wire [0:1] mux_2level_tapbuf_size3_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_60_sram;
wire [0:1] mux_2level_tapbuf_size3_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_61_sram;
wire [0:1] mux_2level_tapbuf_size3_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_62_sram;
wire [0:1] mux_2level_tapbuf_size3_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_63_sram;
wire [0:1] mux_2level_tapbuf_size3_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_64_sram;
wire [0:1] mux_2level_tapbuf_size3_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_65_sram;
wire [0:1] mux_2level_tapbuf_size3_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_66_sram;
wire [0:1] mux_2level_tapbuf_size3_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_67_sram;
wire [0:1] mux_2level_tapbuf_size3_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_68_sram;
wire [0:1] mux_2level_tapbuf_size3_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_69_sram;
wire [0:1] mux_2level_tapbuf_size3_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_70_sram;
wire [0:1] mux_2level_tapbuf_size3_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_71_sram;
wire [0:1] mux_2level_tapbuf_size3_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_72_sram;
wire [0:1] mux_2level_tapbuf_size3_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_73_sram;
wire [0:1] mux_2level_tapbuf_size3_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_74_sram;
wire [0:1] mux_2level_tapbuf_size3_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_75_sram;
wire [0:1] mux_2level_tapbuf_size3_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_76_sram;
wire [0:1] mux_2level_tapbuf_size3_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_77_sram;
wire [0:1] mux_2level_tapbuf_size3_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_78_sram;
wire [0:1] mux_2level_tapbuf_size3_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_79_sram;
wire [0:1] mux_2level_tapbuf_size3_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_80_sram;
wire [0:1] mux_2level_tapbuf_size3_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_81_sram;
wire [0:1] mux_2level_tapbuf_size3_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_82_sram;
wire [0:1] mux_2level_tapbuf_size3_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_83_sram;
wire [0:1] mux_2level_tapbuf_size3_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_84_sram;
wire [0:1] mux_2level_tapbuf_size3_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_85_sram;
wire [0:1] mux_2level_tapbuf_size3_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_86_sram;
wire [0:1] mux_2level_tapbuf_size3_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_87_sram;
wire [0:1] mux_2level_tapbuf_size3_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_88_sram;
wire [0:1] mux_2level_tapbuf_size3_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_89_sram;
wire [0:1] mux_2level_tapbuf_size3_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_8_sram;
wire [0:1] mux_2level_tapbuf_size3_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_90_sram;
wire [0:1] mux_2level_tapbuf_size3_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_91_sram;
wire [0:1] mux_2level_tapbuf_size3_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_92_sram;
wire [0:1] mux_2level_tapbuf_size3_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_93_sram;
wire [0:1] mux_2level_tapbuf_size3_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_94_sram;
wire [0:1] mux_2level_tapbuf_size3_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_95_sram;
wire [0:1] mux_2level_tapbuf_size3_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_96_sram;
wire [0:1] mux_2level_tapbuf_size3_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_97_sram;
wire [0:1] mux_2level_tapbuf_size3_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_98_sram;
wire [0:1] mux_2level_tapbuf_size3_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_99_sram;
wire [0:1] mux_2level_tapbuf_size3_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_9_sram;
wire [0:1] mux_2level_tapbuf_size3_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_144_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_145_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_146_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_147_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_148_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_149_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_150_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_151_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_152_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_153_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_154_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_155_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_156_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_157_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_158_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_159_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_0_sram;
wire [0:5] mux_2level_tapbuf_size8_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_10_sram;
wire [0:5] mux_2level_tapbuf_size8_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_11_sram;
wire [0:5] mux_2level_tapbuf_size8_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_12_sram;
wire [0:5] mux_2level_tapbuf_size8_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_13_sram;
wire [0:5] mux_2level_tapbuf_size8_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_14_sram;
wire [0:5] mux_2level_tapbuf_size8_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_15_sram;
wire [0:5] mux_2level_tapbuf_size8_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_16_sram;
wire [0:5] mux_2level_tapbuf_size8_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_17_sram;
wire [0:5] mux_2level_tapbuf_size8_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_18_sram;
wire [0:5] mux_2level_tapbuf_size8_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_19_sram;
wire [0:5] mux_2level_tapbuf_size8_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_1_sram;
wire [0:5] mux_2level_tapbuf_size8_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_20_sram;
wire [0:5] mux_2level_tapbuf_size8_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_21_sram;
wire [0:5] mux_2level_tapbuf_size8_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_22_sram;
wire [0:5] mux_2level_tapbuf_size8_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_23_sram;
wire [0:5] mux_2level_tapbuf_size8_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_24_sram;
wire [0:5] mux_2level_tapbuf_size8_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_25_sram;
wire [0:5] mux_2level_tapbuf_size8_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_26_sram;
wire [0:5] mux_2level_tapbuf_size8_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_27_sram;
wire [0:5] mux_2level_tapbuf_size8_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_28_sram;
wire [0:5] mux_2level_tapbuf_size8_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_29_sram;
wire [0:5] mux_2level_tapbuf_size8_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_2_sram;
wire [0:5] mux_2level_tapbuf_size8_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_30_sram;
wire [0:5] mux_2level_tapbuf_size8_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_3_sram;
wire [0:5] mux_2level_tapbuf_size8_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_4_sram;
wire [0:5] mux_2level_tapbuf_size8_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_5_sram;
wire [0:5] mux_2level_tapbuf_size8_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_6_sram;
wire [0:5] mux_2level_tapbuf_size8_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_7_sram;
wire [0:5] mux_2level_tapbuf_size8_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_8_sram;
wire [0:5] mux_2level_tapbuf_size8_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size8_9_sram;
wire [0:5] mux_2level_tapbuf_size8_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size8_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size9_0_sram;
wire [0:7] mux_2level_tapbuf_size9_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_1_sram;
wire [0:7] mux_2level_tapbuf_size9_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_2_sram;
wire [0:7] mux_2level_tapbuf_size9_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_3_sram;
wire [0:7] mux_2level_tapbuf_size9_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_4_sram;
wire [0:7] mux_2level_tapbuf_size9_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_5_sram;
wire [0:7] mux_2level_tapbuf_size9_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size9_6_sram;
wire [0:7] mux_2level_tapbuf_size9_6_sram_inv;
wire [0:0] mux_2level_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size9_mem_6_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[1];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[5];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[9];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[13];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[17];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[21];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[25];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[29];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[33];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[37];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[41];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[45];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[49];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[53];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[57];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[61];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[64] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[65];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[68] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[69];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[72] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[73];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[76] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[77];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[80] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[81];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[84] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[85];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[88] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[89];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[92] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[93];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[96] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[97];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[100] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[101];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[104] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[105];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[108] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[109];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[112] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[113];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[116] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[117];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[120] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[121];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[124] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[125];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[128] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[129];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[132] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[133];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[136] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[137];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[140] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[141];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[144] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[145];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[148] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[149];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[152] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[153];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[156] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[157];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[159];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[1];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[5];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[9];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[13];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[17];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[21];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[25];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[29];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[33];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[37];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[41];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[45];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[49];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[53];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[57];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[61];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[64];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[65];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[67];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[68];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[69];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[71];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chany_bottom_in[72];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[73];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[75];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chany_bottom_in[76];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[77];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[79];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chany_bottom_in[80];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[81];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[83];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chany_bottom_in[84];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[85];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[87];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chany_bottom_in[88];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[89];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[91];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chany_bottom_in[92];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[93];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[95];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[96] = chany_bottom_in[96];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[97];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[99];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[100] = chany_bottom_in[100];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[101];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[103];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[104] = chany_bottom_in[104];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[105];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[107];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[108] = chany_bottom_in[108];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[109];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[111];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[112] = chany_bottom_in[112];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[113];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[115];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chany_bottom_in[116];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[117];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[119];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[120] = chany_bottom_in[120];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[121];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[123];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[124] = chany_bottom_in[124];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[125];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[127];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[128] = chany_bottom_in[128];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[129];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[131];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chany_bottom_in[132];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[133];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[135];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[136] = chany_bottom_in[136];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[137];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[139];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[140] = chany_bottom_in[140];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[141];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[143];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[144] = chany_bottom_in[144];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[145];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[147];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[148] = chany_bottom_in[148];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[149];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[151];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chany_bottom_in[152];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[153];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[155];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[156] = chany_bottom_in[156];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[157];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[159];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size11 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[1], chanx_right_in[41], chanx_right_in[81], chanx_right_in[121], chany_bottom_in[2]}),
		.sram(mux_2level_tapbuf_size11_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_0_sram_inv[0:7]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size11 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[2], chanx_right_in[42], chanx_right_in[82], chanx_right_in[122], chany_bottom_in[6]}),
		.sram(mux_2level_tapbuf_size11_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_1_sram_inv[0:7]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size11 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[3], chanx_right_in[43], chanx_right_in[83], chanx_right_in[123], chany_bottom_in[10]}),
		.sram(mux_2level_tapbuf_size11_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_2_sram_inv[0:7]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size11 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[4], chanx_right_in[44], chanx_right_in[84], chanx_right_in[124], chany_bottom_in[14]}),
		.sram(mux_2level_tapbuf_size11_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_3_sram_inv[0:7]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size11 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[5], chanx_right_in[45], chanx_right_in[85], chanx_right_in[125], chany_bottom_in[18]}),
		.sram(mux_2level_tapbuf_size11_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_4_sram_inv[0:7]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size11 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[6], chanx_right_in[46], chanx_right_in[86], chanx_right_in[126], chany_bottom_in[22]}),
		.sram(mux_2level_tapbuf_size11_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_5_sram_inv[0:7]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size11 mux_top_track_52 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[7], chanx_right_in[47], chanx_right_in[87], chanx_right_in[127], chany_bottom_in[26]}),
		.sram(mux_2level_tapbuf_size11_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_6_sram_inv[0:7]),
		.out(chany_top_out[26]));

	mux_2level_tapbuf_size11 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[8], chanx_right_in[48], chanx_right_in[88], chanx_right_in[128], chany_bottom_in[30]}),
		.sram(mux_2level_tapbuf_size11_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_7_sram_inv[0:7]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size11 mux_bottom_track_5 (
		.in({chany_top_in[2], chanx_right_in[38], chanx_right_in[78], chanx_right_in[118], chanx_right_in[158], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size11_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_8_sram_inv[0:7]),
		.out(chany_bottom_out[2]));

	mux_2level_tapbuf_size11_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_0_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_1_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_2_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_3_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_4_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_5_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_6_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_7_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_159_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_8_sram_inv[0:7]));

	mux_2level_tapbuf_size10 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[9], chanx_right_in[49], chanx_right_in[89], chanx_right_in[129], chany_bottom_in[34]}),
		.sram(mux_2level_tapbuf_size10_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_0_sram_inv[0:7]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size10 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[10], chanx_right_in[50], chanx_right_in[90], chanx_right_in[130], chany_bottom_in[38]}),
		.sram(mux_2level_tapbuf_size10_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_1_sram_inv[0:7]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size10 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[11], chanx_right_in[51], chanx_right_in[91], chanx_right_in[131], chany_bottom_in[42]}),
		.sram(mux_2level_tapbuf_size10_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_2_sram_inv[0:7]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size10 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[12], chanx_right_in[52], chanx_right_in[92], chanx_right_in[132], chany_bottom_in[46]}),
		.sram(mux_2level_tapbuf_size10_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_3_sram_inv[0:7]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size10 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[13], chanx_right_in[53], chanx_right_in[93], chanx_right_in[133], chany_bottom_in[50]}),
		.sram(mux_2level_tapbuf_size10_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_4_sram_inv[0:7]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size10 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[14], chanx_right_in[54], chanx_right_in[94], chanx_right_in[134], chany_bottom_in[54]}),
		.sram(mux_2level_tapbuf_size10_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_5_sram_inv[0:7]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size10 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[15], chanx_right_in[55], chanx_right_in[95], chanx_right_in[135], chany_bottom_in[58]}),
		.sram(mux_2level_tapbuf_size10_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_6_sram_inv[0:7]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size10 mux_top_track_124 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[16], chanx_right_in[56], chanx_right_in[96], chanx_right_in[136], chany_bottom_in[62]}),
		.sram(mux_2level_tapbuf_size10_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_7_sram_inv[0:7]),
		.out(chany_top_out[62]));

	mux_2level_tapbuf_size10 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[17], chanx_right_in[57], chanx_right_in[97], chanx_right_in[137], chany_bottom_in[66]}),
		.sram(mux_2level_tapbuf_size10_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_8_sram_inv[0:7]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size10 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[18], chanx_right_in[58], chanx_right_in[98], chanx_right_in[138], chany_bottom_in[70]}),
		.sram(mux_2level_tapbuf_size10_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_9_sram_inv[0:7]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size10 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[19], chanx_right_in[59], chanx_right_in[99], chanx_right_in[139], chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size10_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_10_sram_inv[0:7]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size10 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[20], chanx_right_in[60], chanx_right_in[100], chanx_right_in[140], chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size10_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_11_sram_inv[0:7]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size10 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[21], chanx_right_in[61], chanx_right_in[101], chanx_right_in[141], chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size10_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_12_sram_inv[0:7]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size10 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[22], chanx_right_in[62], chanx_right_in[102], chanx_right_in[142], chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size10_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_13_sram_inv[0:7]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size10 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[23], chanx_right_in[63], chanx_right_in[103], chanx_right_in[143], chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size10_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_14_sram_inv[0:7]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size10 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[24], chanx_right_in[64], chanx_right_in[104], chanx_right_in[144], chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size10_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_15_sram_inv[0:7]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size10 mux_top_track_196 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[25], chanx_right_in[65], chanx_right_in[105], chanx_right_in[145], chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size10_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_16_sram_inv[0:7]),
		.out(chany_top_out[98]));

	mux_2level_tapbuf_size10 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[26], chanx_right_in[66], chanx_right_in[106], chanx_right_in[146], chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size10_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_17_sram_inv[0:7]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size10 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[27], chanx_right_in[67], chanx_right_in[107], chanx_right_in[147], chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size10_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_18_sram_inv[0:7]),
		.out(chany_top_out[106]));

	mux_2level_tapbuf_size10 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[28], chanx_right_in[68], chanx_right_in[108], chanx_right_in[148], chany_bottom_in[110]}),
		.sram(mux_2level_tapbuf_size10_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_19_sram_inv[0:7]),
		.out(chany_top_out[110]));

	mux_2level_tapbuf_size10 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[29], chanx_right_in[69], chanx_right_in[109], chanx_right_in[149], chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size10_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_20_sram_inv[0:7]),
		.out(chany_top_out[114]));

	mux_2level_tapbuf_size10 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[30], chanx_right_in[70], chanx_right_in[110], chanx_right_in[150], chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size10_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_21_sram_inv[0:7]),
		.out(chany_top_out[118]));

	mux_2level_tapbuf_size10 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[31], chanx_right_in[71], chanx_right_in[111], chanx_right_in[151], chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size10_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_22_sram_inv[0:7]),
		.out(chany_top_out[122]));

	mux_2level_tapbuf_size10 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[32], chanx_right_in[72], chanx_right_in[112], chanx_right_in[152], chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size10_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_23_sram_inv[0:7]),
		.out(chany_top_out[126]));

	mux_2level_tapbuf_size10 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[33], chanx_right_in[73], chanx_right_in[113], chanx_right_in[153], chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size10_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_24_sram_inv[0:7]),
		.out(chany_top_out[130]));

	mux_2level_tapbuf_size10 mux_top_track_268 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[34], chanx_right_in[74], chanx_right_in[114], chanx_right_in[154], chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size10_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_25_sram_inv[0:7]),
		.out(chany_top_out[134]));

	mux_2level_tapbuf_size10 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[35], chanx_right_in[75], chanx_right_in[115], chanx_right_in[155], chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size10_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_26_sram_inv[0:7]),
		.out(chany_top_out[138]));

	mux_2level_tapbuf_size10 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[36], chanx_right_in[76], chanx_right_in[116], chanx_right_in[156], chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size10_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_27_sram_inv[0:7]),
		.out(chany_top_out[142]));

	mux_2level_tapbuf_size10 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[37], chanx_right_in[77], chanx_right_in[117], chanx_right_in[157], chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size10_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_28_sram_inv[0:7]),
		.out(chany_top_out[146]));

	mux_2level_tapbuf_size10 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[38], chanx_right_in[78], chanx_right_in[118], chanx_right_in[158], chany_bottom_in[150]}),
		.sram(mux_2level_tapbuf_size10_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_29_sram_inv[0:7]),
		.out(chany_top_out[150]));

	mux_2level_tapbuf_size10 mux_top_track_308 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[39], chanx_right_in[79], chanx_right_in[119], chanx_right_in[159], chany_bottom_in[154]}),
		.sram(mux_2level_tapbuf_size10_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_30_sram_inv[0:7]),
		.out(chany_top_out[154]));

	mux_2level_tapbuf_size10 mux_top_track_316 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[0], chanx_right_in[40], chanx_right_in[80], chanx_right_in[120], chany_bottom_in[158]}),
		.sram(mux_2level_tapbuf_size10_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_31_sram_inv[0:7]),
		.out(chany_top_out[158]));

	mux_2level_tapbuf_size10_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_0_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_1_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_2_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_3_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_4_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_5_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_6_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_7_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_8_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_9_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_10_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_11_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_12_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_13_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_14_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_15_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_16_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_17_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_18_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_19_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_20_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_21_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_22_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_23_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_24_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_25_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_26_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_27_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_28_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_29_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_30_sram_inv[0:7]));

	mux_2level_tapbuf_size10_mem mem_top_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_31_sram_inv[0:7]));

	mux_2level_tapbuf_size3 mux_right_track_0 (
		.in({chany_top_in[159], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[157]}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[2], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[156]}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[6], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[155]}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[10], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[153]}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size3 mux_right_track_8 (
		.in({chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[152]}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size3 mux_right_track_10 (
		.in({chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[151]}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size3 mux_right_track_12 (
		.in({chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[149]}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size3 mux_right_track_14 (
		.in({chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size3 mux_right_track_16 (
		.in({chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[147]}),
		.sram(mux_2level_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size3 mux_right_track_18 (
		.in({chany_top_in[34], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size3 mux_right_track_20 (
		.in({chany_top_in[38], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size3 mux_right_track_22 (
		.in({chany_top_in[42], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[143]}),
		.sram(mux_2level_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size3 mux_right_track_24 (
		.in({chany_top_in[46], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size3 mux_right_track_26 (
		.in({chany_top_in[50], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[140]}),
		.sram(mux_2level_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size3 mux_right_track_28 (
		.in({chany_top_in[54], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[139]}),
		.sram(mux_2level_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size3 mux_right_track_30 (
		.in({chany_top_in[58], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size3 mux_right_track_32 (
		.in({chany_top_in[62], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size3 mux_right_track_34 (
		.in({chany_top_in[66], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[135]}),
		.sram(mux_2level_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size3 mux_right_track_36 (
		.in({chany_top_in[70], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size3 mux_right_track_38 (
		.in({chany_top_in[74], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size3 mux_right_track_40 (
		.in({chany_top_in[78], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[131]}),
		.sram(mux_2level_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size3 mux_right_track_42 (
		.in({chany_top_in[82], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[129]}),
		.sram(mux_2level_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size3 mux_right_track_44 (
		.in({chany_top_in[86], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size3 mux_right_track_46 (
		.in({chany_top_in[90], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[127]}),
		.sram(mux_2level_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size3 mux_right_track_48 (
		.in({chany_top_in[94], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size3 mux_right_track_50 (
		.in({chany_top_in[98], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size3 mux_right_track_52 (
		.in({chany_top_in[102], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[123]}),
		.sram(mux_2level_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size3 mux_right_track_54 (
		.in({chany_top_in[106], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size3 mux_right_track_56 (
		.in({chany_top_in[110], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[120]}),
		.sram(mux_2level_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size3 mux_right_track_58 (
		.in({chany_top_in[114], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[119]}),
		.sram(mux_2level_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size3 mux_right_track_60 (
		.in({chany_top_in[118], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size3 mux_right_track_62 (
		.in({chany_top_in[122], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size3 mux_right_track_64 (
		.in({chany_top_in[126], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[115]}),
		.sram(mux_2level_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size3 mux_right_track_66 (
		.in({chany_top_in[130], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size3 mux_right_track_68 (
		.in({chany_top_in[134], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size3 mux_right_track_70 (
		.in({chany_top_in[138], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[111]}),
		.sram(mux_2level_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_2level_tapbuf_size3 mux_right_track_72 (
		.in({chany_top_in[142], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[109]}),
		.sram(mux_2level_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size3 mux_right_track_74 (
		.in({chany_top_in[146], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[108]}),
		.sram(mux_2level_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size3 mux_right_track_76 (
		.in({chany_top_in[150], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[107]}),
		.sram(mux_2level_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size3 mux_right_track_78 (
		.in({chany_top_in[154], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[105]}),
		.sram(mux_2level_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size3 mux_right_track_80 (
		.in({chany_top_in[158], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size3 mux_right_track_82 (
		.in({chany_top_in[0], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size3 mux_right_track_84 (
		.in({chany_top_in[1], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size3 mux_right_track_86 (
		.in({chany_top_in[3], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size3 mux_right_track_88 (
		.in({chany_top_in[4], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[99]}),
		.sram(mux_2level_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size3 mux_right_track_90 (
		.in({chany_top_in[5], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size3 mux_right_track_92 (
		.in({chany_top_in[7], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size3 mux_right_track_94 (
		.in({chany_top_in[8], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[95]}),
		.sram(mux_2level_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size3 mux_right_track_96 (
		.in({chany_top_in[9], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size3 mux_right_track_98 (
		.in({chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size3 mux_right_track_100 (
		.in({chany_top_in[12], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[91]}),
		.sram(mux_2level_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size3 mux_right_track_102 (
		.in({chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[89]}),
		.sram(mux_2level_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size3 mux_right_track_104 (
		.in({chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size3 mux_right_track_106 (
		.in({chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[87]}),
		.sram(mux_2level_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_2level_tapbuf_size3 mux_right_track_108 (
		.in({chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size3 mux_right_track_110 (
		.in({chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_55_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size3 mux_right_track_112 (
		.in({chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[83]}),
		.sram(mux_2level_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_56_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size3 mux_right_track_114 (
		.in({chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_57_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size3 mux_right_track_116 (
		.in({chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[80]}),
		.sram(mux_2level_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_58_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size3 mux_right_track_118 (
		.in({chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[79]}),
		.sram(mux_2level_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_59_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_2level_tapbuf_size3 mux_right_track_120 (
		.in({chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_60_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size3 mux_right_track_122 (
		.in({chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_61_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size3 mux_right_track_124 (
		.in({chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[75]}),
		.sram(mux_2level_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_62_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_2level_tapbuf_size3 mux_right_track_126 (
		.in({chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_63_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size3 mux_right_track_128 (
		.in({chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[72]}),
		.sram(mux_2level_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_64_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size3 mux_right_track_130 (
		.in({chany_top_in[32], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[71]}),
		.sram(mux_2level_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_65_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size3 mux_right_track_132 (
		.in({chany_top_in[33], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[69]}),
		.sram(mux_2level_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_66_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size3 mux_right_track_134 (
		.in({chany_top_in[35], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[68]}),
		.sram(mux_2level_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_67_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size3 mux_right_track_136 (
		.in({chany_top_in[36], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[67]}),
		.sram(mux_2level_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_68_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size3 mux_right_track_138 (
		.in({chany_top_in[37], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[65]}),
		.sram(mux_2level_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_69_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size3 mux_right_track_140 (
		.in({chany_top_in[39], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[64]}),
		.sram(mux_2level_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_70_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size3 mux_right_track_142 (
		.in({chany_top_in[40], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[63]}),
		.sram(mux_2level_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_71_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_2level_tapbuf_size3 mux_right_track_144 (
		.in({chany_top_in[41], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[61]}),
		.sram(mux_2level_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_72_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size3 mux_right_track_146 (
		.in({chany_top_in[43], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[60]}),
		.sram(mux_2level_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_73_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size3 mux_right_track_148 (
		.in({chany_top_in[44], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[59]}),
		.sram(mux_2level_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_74_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size3 mux_right_track_150 (
		.in({chany_top_in[45], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[57]}),
		.sram(mux_2level_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_75_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size3 mux_right_track_152 (
		.in({chany_top_in[47], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[56]}),
		.sram(mux_2level_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_76_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size3 mux_right_track_154 (
		.in({chany_top_in[48], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[55]}),
		.sram(mux_2level_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_77_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size3 mux_right_track_156 (
		.in({chany_top_in[49], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[53]}),
		.sram(mux_2level_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_78_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size3 mux_right_track_158 (
		.in({chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[52]}),
		.sram(mux_2level_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_79_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_2level_tapbuf_size3 mux_right_track_160 (
		.in({chany_top_in[52], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[51]}),
		.sram(mux_2level_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_80_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size3 mux_right_track_162 (
		.in({chany_top_in[53], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[49]}),
		.sram(mux_2level_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_81_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size3 mux_right_track_164 (
		.in({chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[48]}),
		.sram(mux_2level_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_82_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size3 mux_right_track_166 (
		.in({chany_top_in[56], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[47]}),
		.sram(mux_2level_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_83_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size3 mux_right_track_168 (
		.in({chany_top_in[57], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[45]}),
		.sram(mux_2level_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_84_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size3 mux_right_track_170 (
		.in({chany_top_in[59], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[44]}),
		.sram(mux_2level_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_85_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size3 mux_right_track_172 (
		.in({chany_top_in[60], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[43]}),
		.sram(mux_2level_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size3 mux_right_track_174 (
		.in({chany_top_in[61], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[41]}),
		.sram(mux_2level_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size3 mux_right_track_176 (
		.in({chany_top_in[63], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[40]}),
		.sram(mux_2level_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size3 mux_right_track_178 (
		.in({chany_top_in[64], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[39]}),
		.sram(mux_2level_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_89_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_2level_tapbuf_size3 mux_right_track_180 (
		.in({chany_top_in[65], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[37]}),
		.sram(mux_2level_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_90_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size3 mux_right_track_182 (
		.in({chany_top_in[67], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[36]}),
		.sram(mux_2level_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_91_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size3 mux_right_track_184 (
		.in({chany_top_in[68], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[35]}),
		.sram(mux_2level_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_92_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size3 mux_right_track_186 (
		.in({chany_top_in[69], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[33]}),
		.sram(mux_2level_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_93_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size3 mux_right_track_188 (
		.in({chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[32]}),
		.sram(mux_2level_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_94_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size3 mux_right_track_190 (
		.in({chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[31]}),
		.sram(mux_2level_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_95_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size3 mux_right_track_192 (
		.in({chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[29]}),
		.sram(mux_2level_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_96_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size3 mux_right_track_194 (
		.in({chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[28]}),
		.sram(mux_2level_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_97_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size3 mux_right_track_196 (
		.in({chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[27]}),
		.sram(mux_2level_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_98_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_2level_tapbuf_size3 mux_right_track_198 (
		.in({chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[25]}),
		.sram(mux_2level_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_99_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_2level_tapbuf_size3 mux_right_track_200 (
		.in({chany_top_in[79], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[24]}),
		.sram(mux_2level_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_100_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size3 mux_right_track_202 (
		.in({chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[23]}),
		.sram(mux_2level_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_101_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size3 mux_right_track_204 (
		.in({chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[21]}),
		.sram(mux_2level_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_102_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size3 mux_right_track_206 (
		.in({chany_top_in[83], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[20]}),
		.sram(mux_2level_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_103_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_2level_tapbuf_size3 mux_right_track_208 (
		.in({chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[19]}),
		.sram(mux_2level_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_104_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size3 mux_right_track_210 (
		.in({chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[17]}),
		.sram(mux_2level_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_105_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size3 mux_right_track_212 (
		.in({chany_top_in[87], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[16]}),
		.sram(mux_2level_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_106_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size3 mux_right_track_214 (
		.in({chany_top_in[88], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[15]}),
		.sram(mux_2level_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_107_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_2level_tapbuf_size3 mux_right_track_216 (
		.in({chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[13]}),
		.sram(mux_2level_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_108_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size3 mux_right_track_218 (
		.in({chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[12]}),
		.sram(mux_2level_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_109_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_2level_tapbuf_size3 mux_right_track_220 (
		.in({chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[11]}),
		.sram(mux_2level_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_110_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size3 mux_right_track_222 (
		.in({chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[9]}),
		.sram(mux_2level_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_111_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_2level_tapbuf_size3 mux_right_track_224 (
		.in({chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[8]}),
		.sram(mux_2level_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_112_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size3 mux_right_track_226 (
		.in({chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[7]}),
		.sram(mux_2level_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_113_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size3 mux_right_track_228 (
		.in({chany_top_in[97], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[5]}),
		.sram(mux_2level_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_114_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size3 mux_right_track_230 (
		.in({chany_top_in[99], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[4]}),
		.sram(mux_2level_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_115_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_2level_tapbuf_size3 mux_right_track_232 (
		.in({chany_top_in[100], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[3]}),
		.sram(mux_2level_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_116_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size3 mux_right_track_234 (
		.in({chany_top_in[101], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[1]}),
		.sram(mux_2level_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_117_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size3 mux_right_track_236 (
		.in({chany_top_in[103], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[0]}),
		.sram(mux_2level_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_118_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_2level_tapbuf_size3 mux_right_track_238 (
		.in({chany_top_in[104], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[158]}),
		.sram(mux_2level_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_119_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_2level_tapbuf_size3 mux_right_track_240 (
		.in({chany_top_in[105], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[154]}),
		.sram(mux_2level_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size3 mux_right_track_242 (
		.in({chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[150]}),
		.sram(mux_2level_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size3 mux_right_track_244 (
		.in({chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size3 mux_right_track_246 (
		.in({chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_2level_tapbuf_size3 mux_right_track_248 (
		.in({chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size3 mux_right_track_250 (
		.in({chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_2level_tapbuf_size3 mux_right_track_252 (
		.in({chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size3 mux_right_track_254 (
		.in({chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_2level_tapbuf_size3 mux_right_track_256 (
		.in({chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size3 mux_right_track_258 (
		.in({chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_2level_tapbuf_size3 mux_right_track_260 (
		.in({chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size3 mux_right_track_262 (
		.in({chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[110]}),
		.sram(mux_2level_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_2level_tapbuf_size3 mux_right_track_264 (
		.in({chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size3 mux_right_track_266 (
		.in({chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size3 mux_right_track_268 (
		.in({chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_2level_tapbuf_size3 mux_right_track_270 (
		.in({chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_2level_tapbuf_size3 mux_right_track_272 (
		.in({chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size3 mux_right_track_274 (
		.in({chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_137_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size3 mux_right_track_276 (
		.in({chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_138_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_2level_tapbuf_size3 mux_right_track_278 (
		.in({chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_139_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_2level_tapbuf_size3 mux_right_track_280 (
		.in({chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_140_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size3 mux_right_track_282 (
		.in({chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[70]}),
		.sram(mux_2level_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_141_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size3 mux_right_track_284 (
		.in({chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[66]}),
		.sram(mux_2level_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_142_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size3 mux_right_track_286 (
		.in({chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[62]}),
		.sram(mux_2level_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_143_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_2level_tapbuf_size3 mux_right_track_288 (
		.in({chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[58]}),
		.sram(mux_2level_tapbuf_size3_144_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_144_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size3 mux_right_track_290 (
		.in({chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[54]}),
		.sram(mux_2level_tapbuf_size3_145_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_145_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size3 mux_right_track_292 (
		.in({chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[50]}),
		.sram(mux_2level_tapbuf_size3_146_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_146_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size3 mux_right_track_294 (
		.in({chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[46]}),
		.sram(mux_2level_tapbuf_size3_147_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_147_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_2level_tapbuf_size3 mux_right_track_296 (
		.in({chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[42]}),
		.sram(mux_2level_tapbuf_size3_148_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_148_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size3 mux_right_track_298 (
		.in({chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[38]}),
		.sram(mux_2level_tapbuf_size3_149_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_149_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_2level_tapbuf_size3 mux_right_track_300 (
		.in({chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[34]}),
		.sram(mux_2level_tapbuf_size3_150_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_150_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_2level_tapbuf_size3 mux_right_track_302 (
		.in({chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[30]}),
		.sram(mux_2level_tapbuf_size3_151_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_151_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_2level_tapbuf_size3 mux_right_track_304 (
		.in({chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[26]}),
		.sram(mux_2level_tapbuf_size3_152_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_152_sram_inv[0:1]),
		.out(chanx_right_out[152]));

	mux_2level_tapbuf_size3 mux_right_track_306 (
		.in({chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[22]}),
		.sram(mux_2level_tapbuf_size3_153_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_153_sram_inv[0:1]),
		.out(chanx_right_out[153]));

	mux_2level_tapbuf_size3 mux_right_track_308 (
		.in({chany_top_in[151], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[18]}),
		.sram(mux_2level_tapbuf_size3_154_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_154_sram_inv[0:1]),
		.out(chanx_right_out[154]));

	mux_2level_tapbuf_size3 mux_right_track_310 (
		.in({chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[14]}),
		.sram(mux_2level_tapbuf_size3_155_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_155_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_2level_tapbuf_size3 mux_right_track_312 (
		.in({chany_top_in[153], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[10]}),
		.sram(mux_2level_tapbuf_size3_156_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_156_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_2level_tapbuf_size3 mux_right_track_314 (
		.in({chany_top_in[155], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[6]}),
		.sram(mux_2level_tapbuf_size3_157_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_157_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_2level_tapbuf_size3 mux_right_track_316 (
		.in({chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[2]}),
		.sram(mux_2level_tapbuf_size3_158_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_158_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_2level_tapbuf_size3 mux_right_track_318 (
		.in({chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[159]}),
		.sram(mux_2level_tapbuf_size3_159_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_159_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_2level_tapbuf_size3_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_8_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_9_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_10_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_11_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_12_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_13_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_14_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_15_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_16_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_17_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_18_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_19_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_20_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_21_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_22_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_23_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_24_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_25_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_26_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_27_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_28_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_29_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_30_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_31_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_32_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_33_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_34_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_35_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_36_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_37_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_38_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_39_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_40_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_41_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_42_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_43_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_44_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_45_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_46_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_47_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_48_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_49_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_50_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_51_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_52_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_53_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_54_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_55_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_56_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_57_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_58_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_59_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_60_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_61_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_62_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_63_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_64_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_65_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_66_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_67_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_68_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_69_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_70_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_71_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_72_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_73_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_74_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_75_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_76_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_77_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_78_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_79_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_80_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_81_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_82_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_83_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_84_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_85_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_86_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_87_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_88_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_89_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_90_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_91_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_92_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_93_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_94_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_95_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_96_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_97_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_98_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_99_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_100_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_101_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_102_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_103_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_104_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_105_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_106_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_107_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_108_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_109_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_110_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_111_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_112_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_113_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_114_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_115_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_116_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_117_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_118_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_119_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_120_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_121_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_122_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_123_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_124_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_125_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_126_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_127_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_128_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_129_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_130_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_131_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_132_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_133_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_134_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_135_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_136_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_137_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_138_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_139_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_140_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_141_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_142_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_143_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_144_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_144_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_144_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_144_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_145_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_145_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_145_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_145_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_146_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_146_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_146_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_146_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_147_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_147_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_147_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_147_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_148_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_148_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_148_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_148_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_149_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_149_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_149_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_149_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_150_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_150_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_150_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_302 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_150_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_151_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_151_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_151_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_151_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_152_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_152_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_152_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_152_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_153_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_153_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_153_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_153_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_154_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_154_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_154_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_310 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_154_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_155_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_155_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_155_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_155_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_156_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_156_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_156_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_156_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_157_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_157_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_157_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_157_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_158_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_158_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_158_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_318 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_158_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_159_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_159_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_159_sram_inv[0:1]));

	mux_2level_tapbuf_size9 mux_bottom_track_13 (
		.in({chany_top_in[6], chanx_right_in[37], chanx_right_in[77], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_0_sram_inv[0:7]),
		.out(chany_bottom_out[6]));

	mux_2level_tapbuf_size9 mux_bottom_track_21 (
		.in({chany_top_in[10], chanx_right_in[36], chanx_right_in[76], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_1_sram_inv[0:7]),
		.out(chany_bottom_out[10]));

	mux_2level_tapbuf_size9 mux_bottom_track_29 (
		.in({chany_top_in[14], chanx_right_in[35], chanx_right_in[75], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_2_sram_inv[0:7]),
		.out(chany_bottom_out[14]));

	mux_2level_tapbuf_size9 mux_bottom_track_37 (
		.in({chany_top_in[18], chanx_right_in[34], chanx_right_in[74], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_3_sram_inv[0:7]),
		.out(chany_bottom_out[18]));

	mux_2level_tapbuf_size9 mux_bottom_track_45 (
		.in({chany_top_in[22], chanx_right_in[33], chanx_right_in[73], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_4_sram_inv[0:7]),
		.out(chany_bottom_out[22]));

	mux_2level_tapbuf_size9 mux_bottom_track_53 (
		.in({chany_top_in[26], chanx_right_in[32], chanx_right_in[72], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_5_sram_inv[0:7]),
		.out(chany_bottom_out[26]));

	mux_2level_tapbuf_size9 mux_bottom_track_61 (
		.in({chany_top_in[30], chanx_right_in[31], chanx_right_in[71], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size9_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size9_6_sram_inv[0:7]),
		.out(chany_bottom_out[30]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_0_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_1_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_2_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_37 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_3_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_4_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_5_sram_inv[0:7]));

	mux_2level_tapbuf_size9_mem mem_bottom_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size9_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size9_6_sram_inv[0:7]));

	mux_2level_tapbuf_size8 mux_bottom_track_69 (
		.in({chany_top_in[34], chanx_right_in[30], chanx_right_in[70], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_0_sram_inv[0:5]),
		.out(chany_bottom_out[34]));

	mux_2level_tapbuf_size8 mux_bottom_track_77 (
		.in({chany_top_in[38], chanx_right_in[29], chanx_right_in[69], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_1_sram_inv[0:5]),
		.out(chany_bottom_out[38]));

	mux_2level_tapbuf_size8 mux_bottom_track_85 (
		.in({chany_top_in[42], chanx_right_in[28], chanx_right_in[68], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_2_sram_inv[0:5]),
		.out(chany_bottom_out[42]));

	mux_2level_tapbuf_size8 mux_bottom_track_93 (
		.in({chany_top_in[46], chanx_right_in[27], chanx_right_in[67], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_3_sram_inv[0:5]),
		.out(chany_bottom_out[46]));

	mux_2level_tapbuf_size8 mux_bottom_track_101 (
		.in({chany_top_in[50], chanx_right_in[26], chanx_right_in[66], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_4_sram_inv[0:5]),
		.out(chany_bottom_out[50]));

	mux_2level_tapbuf_size8 mux_bottom_track_109 (
		.in({chany_top_in[54], chanx_right_in[25], chanx_right_in[65], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_5_sram_inv[0:5]),
		.out(chany_bottom_out[54]));

	mux_2level_tapbuf_size8 mux_bottom_track_117 (
		.in({chany_top_in[58], chanx_right_in[24], chanx_right_in[64], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_6_sram_inv[0:5]),
		.out(chany_bottom_out[58]));

	mux_2level_tapbuf_size8 mux_bottom_track_125 (
		.in({chany_top_in[62], chanx_right_in[23], chanx_right_in[63], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_7_sram_inv[0:5]),
		.out(chany_bottom_out[62]));

	mux_2level_tapbuf_size8 mux_bottom_track_133 (
		.in({chany_top_in[66], chanx_right_in[22], chanx_right_in[62], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_8_sram_inv[0:5]),
		.out(chany_bottom_out[66]));

	mux_2level_tapbuf_size8 mux_bottom_track_141 (
		.in({chany_top_in[70], chanx_right_in[21], chanx_right_in[61], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_9_sram_inv[0:5]),
		.out(chany_bottom_out[70]));

	mux_2level_tapbuf_size8 mux_bottom_track_149 (
		.in({chany_top_in[74], chanx_right_in[20], chanx_right_in[60], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_10_sram_inv[0:5]),
		.out(chany_bottom_out[74]));

	mux_2level_tapbuf_size8 mux_bottom_track_157 (
		.in({chany_top_in[78], chanx_right_in[19], chanx_right_in[59], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_11_sram_inv[0:5]),
		.out(chany_bottom_out[78]));

	mux_2level_tapbuf_size8 mux_bottom_track_165 (
		.in({chany_top_in[82], chanx_right_in[18], chanx_right_in[58], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_12_sram_inv[0:5]),
		.out(chany_bottom_out[82]));

	mux_2level_tapbuf_size8 mux_bottom_track_173 (
		.in({chany_top_in[86], chanx_right_in[17], chanx_right_in[57], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_13_sram_inv[0:5]),
		.out(chany_bottom_out[86]));

	mux_2level_tapbuf_size8 mux_bottom_track_181 (
		.in({chany_top_in[90], chanx_right_in[16], chanx_right_in[56], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_14_sram_inv[0:5]),
		.out(chany_bottom_out[90]));

	mux_2level_tapbuf_size8 mux_bottom_track_189 (
		.in({chany_top_in[94], chanx_right_in[15], chanx_right_in[55], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_15_sram_inv[0:5]),
		.out(chany_bottom_out[94]));

	mux_2level_tapbuf_size8 mux_bottom_track_197 (
		.in({chany_top_in[98], chanx_right_in[14], chanx_right_in[54], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_16_sram_inv[0:5]),
		.out(chany_bottom_out[98]));

	mux_2level_tapbuf_size8 mux_bottom_track_205 (
		.in({chany_top_in[102], chanx_right_in[13], chanx_right_in[53], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_17_sram_inv[0:5]),
		.out(chany_bottom_out[102]));

	mux_2level_tapbuf_size8 mux_bottom_track_213 (
		.in({chany_top_in[106], chanx_right_in[12], chanx_right_in[52], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_18_sram_inv[0:5]),
		.out(chany_bottom_out[106]));

	mux_2level_tapbuf_size8 mux_bottom_track_221 (
		.in({chany_top_in[110], chanx_right_in[11], chanx_right_in[51], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_19_sram_inv[0:5]),
		.out(chany_bottom_out[110]));

	mux_2level_tapbuf_size8 mux_bottom_track_229 (
		.in({chany_top_in[114], chanx_right_in[10], chanx_right_in[50], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_20_sram_inv[0:5]),
		.out(chany_bottom_out[114]));

	mux_2level_tapbuf_size8 mux_bottom_track_237 (
		.in({chany_top_in[118], chanx_right_in[9], chanx_right_in[49], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_21_sram_inv[0:5]),
		.out(chany_bottom_out[118]));

	mux_2level_tapbuf_size8 mux_bottom_track_245 (
		.in({chany_top_in[122], chanx_right_in[8], chanx_right_in[48], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_22_sram_inv[0:5]),
		.out(chany_bottom_out[122]));

	mux_2level_tapbuf_size8 mux_bottom_track_253 (
		.in({chany_top_in[126], chanx_right_in[7], chanx_right_in[47], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_23_sram_inv[0:5]),
		.out(chany_bottom_out[126]));

	mux_2level_tapbuf_size8 mux_bottom_track_261 (
		.in({chany_top_in[130], chanx_right_in[6], chanx_right_in[46], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_24_sram_inv[0:5]),
		.out(chany_bottom_out[130]));

	mux_2level_tapbuf_size8 mux_bottom_track_269 (
		.in({chany_top_in[134], chanx_right_in[5], chanx_right_in[45], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_25_sram_inv[0:5]),
		.out(chany_bottom_out[134]));

	mux_2level_tapbuf_size8 mux_bottom_track_277 (
		.in({chany_top_in[138], chanx_right_in[4], chanx_right_in[44], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_26_sram_inv[0:5]),
		.out(chany_bottom_out[138]));

	mux_2level_tapbuf_size8 mux_bottom_track_285 (
		.in({chany_top_in[142], chanx_right_in[3], chanx_right_in[43], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_27_sram_inv[0:5]),
		.out(chany_bottom_out[142]));

	mux_2level_tapbuf_size8 mux_bottom_track_293 (
		.in({chany_top_in[146], chanx_right_in[2], chanx_right_in[42], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_28_sram_inv[0:5]),
		.out(chany_bottom_out[146]));

	mux_2level_tapbuf_size8 mux_bottom_track_301 (
		.in({chany_top_in[150], chanx_right_in[1], chanx_right_in[41], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_29_sram_inv[0:5]),
		.out(chany_bottom_out[150]));

	mux_2level_tapbuf_size8 mux_bottom_track_309 (
		.in({chany_top_in[154], chanx_right_in[0], chanx_right_in[40], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size8_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size8_30_sram_inv[0:5]),
		.out(chany_bottom_out[154]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_0_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_77 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_1_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_2_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_3_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_101 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_4_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_109 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_5_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_117 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_6_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_125 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_7_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_133 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_8_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_141 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_9_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_149 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_10_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_157 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_11_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_165 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_12_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_173 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_13_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_181 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_14_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_189 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_15_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_197 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_16_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_205 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_17_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_213 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_18_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_221 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_19_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_229 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_20_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_237 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_21_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_245 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_22_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_253 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_23_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_261 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_24_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_269 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_25_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_277 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_26_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_285 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_27_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_293 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_28_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_301 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_29_sram_inv[0:5]));

	mux_2level_tapbuf_size8_mem mem_bottom_track_309 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size8_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size8_30_sram_inv[0:5]));

	mux_2level_tapbuf_size7 mux_bottom_track_317 (
		.in({chany_top_in[158], chanx_right_in[39], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_bottom_out[158]));

	mux_2level_tapbuf_size7_mem mem_bottom_track_317 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

endmodule
// ----- END Verilog module for sb_0__2_ -----

//----- Default net type -----
`default_nettype wire



