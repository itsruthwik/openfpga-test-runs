//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Sep 25 15:37:36 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__4_ -----
module sb_0__4_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:216] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:216] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:216] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:216] chany_top_out;
//----- OUTPUT PORTS -----
output [0:216] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:216] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_100_sram;
wire [0:1] mux_2level_tapbuf_size2_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_101_sram;
wire [0:1] mux_2level_tapbuf_size2_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_102_sram;
wire [0:1] mux_2level_tapbuf_size2_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_103_sram;
wire [0:1] mux_2level_tapbuf_size2_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_104_sram;
wire [0:1] mux_2level_tapbuf_size2_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_105_sram;
wire [0:1] mux_2level_tapbuf_size2_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_106_sram;
wire [0:1] mux_2level_tapbuf_size2_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_107_sram;
wire [0:1] mux_2level_tapbuf_size2_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_108_sram;
wire [0:1] mux_2level_tapbuf_size2_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_109_sram;
wire [0:1] mux_2level_tapbuf_size2_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_110_sram;
wire [0:1] mux_2level_tapbuf_size2_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_111_sram;
wire [0:1] mux_2level_tapbuf_size2_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_60_sram;
wire [0:1] mux_2level_tapbuf_size2_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_61_sram;
wire [0:1] mux_2level_tapbuf_size2_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_62_sram;
wire [0:1] mux_2level_tapbuf_size2_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_63_sram;
wire [0:1] mux_2level_tapbuf_size2_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_64_sram;
wire [0:1] mux_2level_tapbuf_size2_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_65_sram;
wire [0:1] mux_2level_tapbuf_size2_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_66_sram;
wire [0:1] mux_2level_tapbuf_size2_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_67_sram;
wire [0:1] mux_2level_tapbuf_size2_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_68_sram;
wire [0:1] mux_2level_tapbuf_size2_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_69_sram;
wire [0:1] mux_2level_tapbuf_size2_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_70_sram;
wire [0:1] mux_2level_tapbuf_size2_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_71_sram;
wire [0:1] mux_2level_tapbuf_size2_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_72_sram;
wire [0:1] mux_2level_tapbuf_size2_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_73_sram;
wire [0:1] mux_2level_tapbuf_size2_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_74_sram;
wire [0:1] mux_2level_tapbuf_size2_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_75_sram;
wire [0:1] mux_2level_tapbuf_size2_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_76_sram;
wire [0:1] mux_2level_tapbuf_size2_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_77_sram;
wire [0:1] mux_2level_tapbuf_size2_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_78_sram;
wire [0:1] mux_2level_tapbuf_size2_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_79_sram;
wire [0:1] mux_2level_tapbuf_size2_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_80_sram;
wire [0:1] mux_2level_tapbuf_size2_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_81_sram;
wire [0:1] mux_2level_tapbuf_size2_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_82_sram;
wire [0:1] mux_2level_tapbuf_size2_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_83_sram;
wire [0:1] mux_2level_tapbuf_size2_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_84_sram;
wire [0:1] mux_2level_tapbuf_size2_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_85_sram;
wire [0:1] mux_2level_tapbuf_size2_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_86_sram;
wire [0:1] mux_2level_tapbuf_size2_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_87_sram;
wire [0:1] mux_2level_tapbuf_size2_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_88_sram;
wire [0:1] mux_2level_tapbuf_size2_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_89_sram;
wire [0:1] mux_2level_tapbuf_size2_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_90_sram;
wire [0:1] mux_2level_tapbuf_size2_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_91_sram;
wire [0:1] mux_2level_tapbuf_size2_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_92_sram;
wire [0:1] mux_2level_tapbuf_size2_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_93_sram;
wire [0:1] mux_2level_tapbuf_size2_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_94_sram;
wire [0:1] mux_2level_tapbuf_size2_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_95_sram;
wire [0:1] mux_2level_tapbuf_size2_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_96_sram;
wire [0:1] mux_2level_tapbuf_size2_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_97_sram;
wire [0:1] mux_2level_tapbuf_size2_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_98_sram;
wire [0:1] mux_2level_tapbuf_size2_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_99_sram;
wire [0:1] mux_2level_tapbuf_size2_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_10_sram;
wire [0:1] mux_2level_tapbuf_size3_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_11_sram;
wire [0:1] mux_2level_tapbuf_size3_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_12_sram;
wire [0:1] mux_2level_tapbuf_size3_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_13_sram;
wire [0:1] mux_2level_tapbuf_size3_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_14_sram;
wire [0:1] mux_2level_tapbuf_size3_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_15_sram;
wire [0:1] mux_2level_tapbuf_size3_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_16_sram;
wire [0:1] mux_2level_tapbuf_size3_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_17_sram;
wire [0:1] mux_2level_tapbuf_size3_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_18_sram;
wire [0:1] mux_2level_tapbuf_size3_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_19_sram;
wire [0:1] mux_2level_tapbuf_size3_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_20_sram;
wire [0:1] mux_2level_tapbuf_size3_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_21_sram;
wire [0:1] mux_2level_tapbuf_size3_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_22_sram;
wire [0:1] mux_2level_tapbuf_size3_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_23_sram;
wire [0:1] mux_2level_tapbuf_size3_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_24_sram;
wire [0:1] mux_2level_tapbuf_size3_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_25_sram;
wire [0:1] mux_2level_tapbuf_size3_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_26_sram;
wire [0:1] mux_2level_tapbuf_size3_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_27_sram;
wire [0:1] mux_2level_tapbuf_size3_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_28_sram;
wire [0:1] mux_2level_tapbuf_size3_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_29_sram;
wire [0:1] mux_2level_tapbuf_size3_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_30_sram;
wire [0:1] mux_2level_tapbuf_size3_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_31_sram;
wire [0:1] mux_2level_tapbuf_size3_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_32_sram;
wire [0:1] mux_2level_tapbuf_size3_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_33_sram;
wire [0:1] mux_2level_tapbuf_size3_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_34_sram;
wire [0:1] mux_2level_tapbuf_size3_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_35_sram;
wire [0:1] mux_2level_tapbuf_size3_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_36_sram;
wire [0:1] mux_2level_tapbuf_size3_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_37_sram;
wire [0:1] mux_2level_tapbuf_size3_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_38_sram;
wire [0:1] mux_2level_tapbuf_size3_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_39_sram;
wire [0:1] mux_2level_tapbuf_size3_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_40_sram;
wire [0:1] mux_2level_tapbuf_size3_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_41_sram;
wire [0:1] mux_2level_tapbuf_size3_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_42_sram;
wire [0:1] mux_2level_tapbuf_size3_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_43_sram;
wire [0:1] mux_2level_tapbuf_size3_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_44_sram;
wire [0:1] mux_2level_tapbuf_size3_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_45_sram;
wire [0:1] mux_2level_tapbuf_size3_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_46_sram;
wire [0:1] mux_2level_tapbuf_size3_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_47_sram;
wire [0:1] mux_2level_tapbuf_size3_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_48_sram;
wire [0:1] mux_2level_tapbuf_size3_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_49_sram;
wire [0:1] mux_2level_tapbuf_size3_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_50_sram;
wire [0:1] mux_2level_tapbuf_size3_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_51_sram;
wire [0:1] mux_2level_tapbuf_size3_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_52_sram;
wire [0:1] mux_2level_tapbuf_size3_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_53_sram;
wire [0:1] mux_2level_tapbuf_size3_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_54_sram;
wire [0:1] mux_2level_tapbuf_size3_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_55_sram;
wire [0:1] mux_2level_tapbuf_size3_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_56_sram;
wire [0:1] mux_2level_tapbuf_size3_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_57_sram;
wire [0:1] mux_2level_tapbuf_size3_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_58_sram;
wire [0:1] mux_2level_tapbuf_size3_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_59_sram;
wire [0:1] mux_2level_tapbuf_size3_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_60_sram;
wire [0:1] mux_2level_tapbuf_size3_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_61_sram;
wire [0:1] mux_2level_tapbuf_size3_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_62_sram;
wire [0:1] mux_2level_tapbuf_size3_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_63_sram;
wire [0:1] mux_2level_tapbuf_size3_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_64_sram;
wire [0:1] mux_2level_tapbuf_size3_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_65_sram;
wire [0:1] mux_2level_tapbuf_size3_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_66_sram;
wire [0:1] mux_2level_tapbuf_size3_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_67_sram;
wire [0:1] mux_2level_tapbuf_size3_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_68_sram;
wire [0:1] mux_2level_tapbuf_size3_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_69_sram;
wire [0:1] mux_2level_tapbuf_size3_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_70_sram;
wire [0:1] mux_2level_tapbuf_size3_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_71_sram;
wire [0:1] mux_2level_tapbuf_size3_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_72_sram;
wire [0:1] mux_2level_tapbuf_size3_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_73_sram;
wire [0:1] mux_2level_tapbuf_size3_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_74_sram;
wire [0:1] mux_2level_tapbuf_size3_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_75_sram;
wire [0:1] mux_2level_tapbuf_size3_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_76_sram;
wire [0:1] mux_2level_tapbuf_size3_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_77_sram;
wire [0:1] mux_2level_tapbuf_size3_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_78_sram;
wire [0:1] mux_2level_tapbuf_size3_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_79_sram;
wire [0:1] mux_2level_tapbuf_size3_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_80_sram;
wire [0:1] mux_2level_tapbuf_size3_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_81_sram;
wire [0:1] mux_2level_tapbuf_size3_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_82_sram;
wire [0:1] mux_2level_tapbuf_size3_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_83_sram;
wire [0:1] mux_2level_tapbuf_size3_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_84_sram;
wire [0:1] mux_2level_tapbuf_size3_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_85_sram;
wire [0:1] mux_2level_tapbuf_size3_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_86_sram;
wire [0:1] mux_2level_tapbuf_size3_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_87_sram;
wire [0:1] mux_2level_tapbuf_size3_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_88_sram;
wire [0:1] mux_2level_tapbuf_size3_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_8_sram;
wire [0:1] mux_2level_tapbuf_size3_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_9_sram;
wire [0:1] mux_2level_tapbuf_size3_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size4_0_sram;
wire [0:5] mux_2level_tapbuf_size4_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_10_sram;
wire [0:5] mux_2level_tapbuf_size4_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_11_sram;
wire [0:5] mux_2level_tapbuf_size4_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_12_sram;
wire [0:5] mux_2level_tapbuf_size4_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_13_sram;
wire [0:5] mux_2level_tapbuf_size4_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_14_sram;
wire [0:5] mux_2level_tapbuf_size4_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_15_sram;
wire [0:5] mux_2level_tapbuf_size4_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_16_sram;
wire [0:5] mux_2level_tapbuf_size4_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_17_sram;
wire [0:5] mux_2level_tapbuf_size4_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_18_sram;
wire [0:5] mux_2level_tapbuf_size4_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_19_sram;
wire [0:5] mux_2level_tapbuf_size4_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_1_sram;
wire [0:5] mux_2level_tapbuf_size4_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_20_sram;
wire [0:5] mux_2level_tapbuf_size4_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_21_sram;
wire [0:5] mux_2level_tapbuf_size4_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_22_sram;
wire [0:5] mux_2level_tapbuf_size4_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_23_sram;
wire [0:5] mux_2level_tapbuf_size4_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_2_sram;
wire [0:5] mux_2level_tapbuf_size4_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_3_sram;
wire [0:5] mux_2level_tapbuf_size4_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_4_sram;
wire [0:5] mux_2level_tapbuf_size4_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_5_sram;
wire [0:5] mux_2level_tapbuf_size4_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_6_sram;
wire [0:5] mux_2level_tapbuf_size4_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_7_sram;
wire [0:5] mux_2level_tapbuf_size4_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_8_sram;
wire [0:5] mux_2level_tapbuf_size4_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size4_9_sram;
wire [0:5] mux_2level_tapbuf_size4_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size4_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size5_0_sram;
wire [0:5] mux_2level_tapbuf_size5_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_10_sram;
wire [0:5] mux_2level_tapbuf_size5_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_11_sram;
wire [0:5] mux_2level_tapbuf_size5_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_12_sram;
wire [0:5] mux_2level_tapbuf_size5_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_13_sram;
wire [0:5] mux_2level_tapbuf_size5_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_14_sram;
wire [0:5] mux_2level_tapbuf_size5_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_15_sram;
wire [0:5] mux_2level_tapbuf_size5_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_16_sram;
wire [0:5] mux_2level_tapbuf_size5_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_17_sram;
wire [0:5] mux_2level_tapbuf_size5_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_18_sram;
wire [0:5] mux_2level_tapbuf_size5_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_19_sram;
wire [0:5] mux_2level_tapbuf_size5_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_1_sram;
wire [0:5] mux_2level_tapbuf_size5_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_20_sram;
wire [0:5] mux_2level_tapbuf_size5_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_21_sram;
wire [0:5] mux_2level_tapbuf_size5_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_22_sram;
wire [0:5] mux_2level_tapbuf_size5_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_23_sram;
wire [0:5] mux_2level_tapbuf_size5_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_24_sram;
wire [0:5] mux_2level_tapbuf_size5_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_25_sram;
wire [0:5] mux_2level_tapbuf_size5_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_26_sram;
wire [0:5] mux_2level_tapbuf_size5_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_27_sram;
wire [0:5] mux_2level_tapbuf_size5_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_28_sram;
wire [0:5] mux_2level_tapbuf_size5_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_29_sram;
wire [0:5] mux_2level_tapbuf_size5_29_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_2_sram;
wire [0:5] mux_2level_tapbuf_size5_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_30_sram;
wire [0:5] mux_2level_tapbuf_size5_30_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_31_sram;
wire [0:5] mux_2level_tapbuf_size5_31_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_32_sram;
wire [0:5] mux_2level_tapbuf_size5_32_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_33_sram;
wire [0:5] mux_2level_tapbuf_size5_33_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_34_sram;
wire [0:5] mux_2level_tapbuf_size5_34_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_35_sram;
wire [0:5] mux_2level_tapbuf_size5_35_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_36_sram;
wire [0:5] mux_2level_tapbuf_size5_36_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_37_sram;
wire [0:5] mux_2level_tapbuf_size5_37_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_38_sram;
wire [0:5] mux_2level_tapbuf_size5_38_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_39_sram;
wire [0:5] mux_2level_tapbuf_size5_39_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_3_sram;
wire [0:5] mux_2level_tapbuf_size5_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_40_sram;
wire [0:5] mux_2level_tapbuf_size5_40_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_41_sram;
wire [0:5] mux_2level_tapbuf_size5_41_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_42_sram;
wire [0:5] mux_2level_tapbuf_size5_42_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_43_sram;
wire [0:5] mux_2level_tapbuf_size5_43_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_44_sram;
wire [0:5] mux_2level_tapbuf_size5_44_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_45_sram;
wire [0:5] mux_2level_tapbuf_size5_45_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_46_sram;
wire [0:5] mux_2level_tapbuf_size5_46_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_47_sram;
wire [0:5] mux_2level_tapbuf_size5_47_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_48_sram;
wire [0:5] mux_2level_tapbuf_size5_48_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_49_sram;
wire [0:5] mux_2level_tapbuf_size5_49_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_4_sram;
wire [0:5] mux_2level_tapbuf_size5_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_50_sram;
wire [0:5] mux_2level_tapbuf_size5_50_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_51_sram;
wire [0:5] mux_2level_tapbuf_size5_51_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_52_sram;
wire [0:5] mux_2level_tapbuf_size5_52_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_53_sram;
wire [0:5] mux_2level_tapbuf_size5_53_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_54_sram;
wire [0:5] mux_2level_tapbuf_size5_54_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_55_sram;
wire [0:5] mux_2level_tapbuf_size5_55_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_56_sram;
wire [0:5] mux_2level_tapbuf_size5_56_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_57_sram;
wire [0:5] mux_2level_tapbuf_size5_57_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_58_sram;
wire [0:5] mux_2level_tapbuf_size5_58_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_59_sram;
wire [0:5] mux_2level_tapbuf_size5_59_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_5_sram;
wire [0:5] mux_2level_tapbuf_size5_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_60_sram;
wire [0:5] mux_2level_tapbuf_size5_60_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_61_sram;
wire [0:5] mux_2level_tapbuf_size5_61_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_62_sram;
wire [0:5] mux_2level_tapbuf_size5_62_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_63_sram;
wire [0:5] mux_2level_tapbuf_size5_63_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_64_sram;
wire [0:5] mux_2level_tapbuf_size5_64_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_65_sram;
wire [0:5] mux_2level_tapbuf_size5_65_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_6_sram;
wire [0:5] mux_2level_tapbuf_size5_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_7_sram;
wire [0:5] mux_2level_tapbuf_size5_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_8_sram;
wire [0:5] mux_2level_tapbuf_size5_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size5_9_sram;
wire [0:5] mux_2level_tapbuf_size5_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size5_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size6_0_sram;
wire [0:5] mux_2level_tapbuf_size6_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_10_sram;
wire [0:5] mux_2level_tapbuf_size6_10_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_11_sram;
wire [0:5] mux_2level_tapbuf_size6_11_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_12_sram;
wire [0:5] mux_2level_tapbuf_size6_12_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_13_sram;
wire [0:5] mux_2level_tapbuf_size6_13_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_14_sram;
wire [0:5] mux_2level_tapbuf_size6_14_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_15_sram;
wire [0:5] mux_2level_tapbuf_size6_15_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_16_sram;
wire [0:5] mux_2level_tapbuf_size6_16_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_17_sram;
wire [0:5] mux_2level_tapbuf_size6_17_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_18_sram;
wire [0:5] mux_2level_tapbuf_size6_18_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_19_sram;
wire [0:5] mux_2level_tapbuf_size6_19_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_1_sram;
wire [0:5] mux_2level_tapbuf_size6_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_20_sram;
wire [0:5] mux_2level_tapbuf_size6_20_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_21_sram;
wire [0:5] mux_2level_tapbuf_size6_21_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_22_sram;
wire [0:5] mux_2level_tapbuf_size6_22_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_23_sram;
wire [0:5] mux_2level_tapbuf_size6_23_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_24_sram;
wire [0:5] mux_2level_tapbuf_size6_24_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_25_sram;
wire [0:5] mux_2level_tapbuf_size6_25_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_26_sram;
wire [0:5] mux_2level_tapbuf_size6_26_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_27_sram;
wire [0:5] mux_2level_tapbuf_size6_27_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_28_sram;
wire [0:5] mux_2level_tapbuf_size6_28_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_2_sram;
wire [0:5] mux_2level_tapbuf_size6_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_3_sram;
wire [0:5] mux_2level_tapbuf_size6_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_4_sram;
wire [0:5] mux_2level_tapbuf_size6_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_5_sram;
wire [0:5] mux_2level_tapbuf_size6_5_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_6_sram;
wire [0:5] mux_2level_tapbuf_size6_6_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_7_sram;
wire [0:5] mux_2level_tapbuf_size6_7_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_8_sram;
wire [0:5] mux_2level_tapbuf_size6_8_sram_inv;
wire [0:5] mux_2level_tapbuf_size6_9_sram;
wire [0:5] mux_2level_tapbuf_size6_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size6_mem_9_ccff_tail;
wire [0:5] mux_2level_tapbuf_size7_0_sram;
wire [0:5] mux_2level_tapbuf_size7_0_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_1_sram;
wire [0:5] mux_2level_tapbuf_size7_1_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_2_sram;
wire [0:5] mux_2level_tapbuf_size7_2_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_3_sram;
wire [0:5] mux_2level_tapbuf_size7_3_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_4_sram;
wire [0:5] mux_2level_tapbuf_size7_4_sram_inv;
wire [0:5] mux_2level_tapbuf_size7_5_sram;
wire [0:5] mux_2level_tapbuf_size7_5_sram_inv;
wire [0:0] mux_2level_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size7_mem_5_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[193] = chany_top_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[194] = chany_top_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[195] = chany_top_in[194];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[197] = chany_top_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[198] = chany_top_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[199] = chany_top_in[198];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[201] = chany_top_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[202] = chany_top_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[203] = chany_top_in[202];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[205] = chany_top_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[206] = chany_top_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[207] = chany_top_in[206];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[209] = chany_top_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[210] = chany_top_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[211] = chany_top_in[210];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[213] = chany_top_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[214] = chany_top_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[215] = chany_top_in[214];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 24 -----
	assign chanx_right_out[216] = right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_[0];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[193] = chany_bottom_in[192];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[194] = chany_bottom_in[193];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[195] = chany_bottom_in[194];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chany_bottom_in[196];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[198] = chany_bottom_in[197];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[199] = chany_bottom_in[198];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[201] = chany_bottom_in[200];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[202] = chany_bottom_in[201];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[203] = chany_bottom_in[202];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[205] = chany_bottom_in[204];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chany_bottom_in[205];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[207] = chany_bottom_in[206];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[209] = chany_bottom_in[208];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[210] = chany_bottom_in[209];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[211] = chany_bottom_in[210];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[213] = chany_bottom_in[212];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[214] = chany_bottom_in[213];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chany_bottom_in[214];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size7 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[1], chanx_right_in[56], chanx_right_in[111], chanx_right_in[166]}),
		.sram(mux_2level_tapbuf_size7_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_0_sram_inv[0:5]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size7 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[2], chanx_right_in[57], chanx_right_in[112], chanx_right_in[167]}),
		.sram(mux_2level_tapbuf_size7_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_1_sram_inv[0:5]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size7 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[3], chanx_right_in[58], chanx_right_in[113], chanx_right_in[168]}),
		.sram(mux_2level_tapbuf_size7_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_2_sram_inv[0:5]),
		.out(chany_top_out[8]));

	mux_2level_tapbuf_size7 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[10], chanx_right_in[65], chanx_right_in[120], chanx_right_in[175]}),
		.sram(mux_2level_tapbuf_size7_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_3_sram_inv[0:5]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size7 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[11], chanx_right_in[66], chanx_right_in[121], chanx_right_in[176]}),
		.sram(mux_2level_tapbuf_size7_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_4_sram_inv[0:5]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size7 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[12], chanx_right_in[67], chanx_right_in[122], chanx_right_in[177]}),
		.sram(mux_2level_tapbuf_size7_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size7_5_sram_inv[0:5]),
		.out(chany_top_out[44]));

	mux_2level_tapbuf_size7_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_0_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_1_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_2_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_3_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_4_sram_inv[0:5]));

	mux_2level_tapbuf_size7_mem mem_top_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size7_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size7_5_sram_inv[0:5]));

	mux_2level_tapbuf_size6 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[4], chanx_right_in[59], chanx_right_in[114], chanx_right_in[169]}),
		.sram(mux_2level_tapbuf_size6_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_0_sram_inv[0:5]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size6 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[5], chanx_right_in[60], chanx_right_in[115], chanx_right_in[170]}),
		.sram(mux_2level_tapbuf_size6_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_1_sram_inv[0:5]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size6 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[6], chanx_right_in[61], chanx_right_in[116], chanx_right_in[171]}),
		.sram(mux_2level_tapbuf_size6_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_2_sram_inv[0:5]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size6 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[7], chanx_right_in[62], chanx_right_in[117], chanx_right_in[172]}),
		.sram(mux_2level_tapbuf_size6_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_3_sram_inv[0:5]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size6 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[8], chanx_right_in[63], chanx_right_in[118], chanx_right_in[173]}),
		.sram(mux_2level_tapbuf_size6_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_4_sram_inv[0:5]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size6 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[9], chanx_right_in[64], chanx_right_in[119], chanx_right_in[174]}),
		.sram(mux_2level_tapbuf_size6_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_5_sram_inv[0:5]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size6 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[13], chanx_right_in[68], chanx_right_in[123], chanx_right_in[178]}),
		.sram(mux_2level_tapbuf_size6_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_6_sram_inv[0:5]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[19], chanx_right_in[74], chanx_right_in[129], chanx_right_in[184]}),
		.sram(mux_2level_tapbuf_size6_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_7_sram_inv[0:5]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size6 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[20], chanx_right_in[75], chanx_right_in[130], chanx_right_in[185]}),
		.sram(mux_2level_tapbuf_size6_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_8_sram_inv[0:5]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size6 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[21], chanx_right_in[76], chanx_right_in[131], chanx_right_in[186]}),
		.sram(mux_2level_tapbuf_size6_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_9_sram_inv[0:5]),
		.out(chany_top_out[80]));

	mux_2level_tapbuf_size6 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[22], chanx_right_in[77], chanx_right_in[132], chanx_right_in[187]}),
		.sram(mux_2level_tapbuf_size6_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_10_sram_inv[0:5]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size6 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[28], chanx_right_in[83], chanx_right_in[138], chanx_right_in[193]}),
		.sram(mux_2level_tapbuf_size6_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_11_sram_inv[0:5]),
		.out(chany_top_out[108]));

	mux_2level_tapbuf_size6 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[29], chanx_right_in[84], chanx_right_in[139], chanx_right_in[194]}),
		.sram(mux_2level_tapbuf_size6_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_12_sram_inv[0:5]),
		.out(chany_top_out[112]));

	mux_2level_tapbuf_size6 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[30], chanx_right_in[85], chanx_right_in[140], chanx_right_in[195]}),
		.sram(mux_2level_tapbuf_size6_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_13_sram_inv[0:5]),
		.out(chany_top_out[116]));

	mux_2level_tapbuf_size6 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[31], chanx_right_in[86], chanx_right_in[141], chanx_right_in[196]}),
		.sram(mux_2level_tapbuf_size6_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_14_sram_inv[0:5]),
		.out(chany_top_out[120]));

	mux_2level_tapbuf_size6 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[37], chanx_right_in[92], chanx_right_in[147], chanx_right_in[202]}),
		.sram(mux_2level_tapbuf_size6_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_15_sram_inv[0:5]),
		.out(chany_top_out[144]));

	mux_2level_tapbuf_size6 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[38], chanx_right_in[93], chanx_right_in[148], chanx_right_in[203]}),
		.sram(mux_2level_tapbuf_size6_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_16_sram_inv[0:5]),
		.out(chany_top_out[148]));

	mux_2level_tapbuf_size6 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[39], chanx_right_in[94], chanx_right_in[149], chanx_right_in[204]}),
		.sram(mux_2level_tapbuf_size6_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_17_sram_inv[0:5]),
		.out(chany_top_out[152]));

	mux_2level_tapbuf_size6 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[40], chanx_right_in[95], chanx_right_in[150], chanx_right_in[205]}),
		.sram(mux_2level_tapbuf_size6_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_18_sram_inv[0:5]),
		.out(chany_top_out[156]));

	mux_2level_tapbuf_size6 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[46], chanx_right_in[101], chanx_right_in[156], chanx_right_in[211]}),
		.sram(mux_2level_tapbuf_size6_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_19_sram_inv[0:5]),
		.out(chany_top_out[180]));

	mux_2level_tapbuf_size6 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[47], chanx_right_in[102], chanx_right_in[157], chanx_right_in[212]}),
		.sram(mux_2level_tapbuf_size6_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_20_sram_inv[0:5]),
		.out(chany_top_out[184]));

	mux_2level_tapbuf_size6 mux_top_track_376 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[48], chanx_right_in[103], chanx_right_in[158], chanx_right_in[213]}),
		.sram(mux_2level_tapbuf_size6_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_21_sram_inv[0:5]),
		.out(chany_top_out[188]));

	mux_2level_tapbuf_size6 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[49], chanx_right_in[104], chanx_right_in[159], chanx_right_in[214]}),
		.sram(mux_2level_tapbuf_size6_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_22_sram_inv[0:5]),
		.out(chany_top_out[192]));

	mux_2level_tapbuf_size6 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, chanx_right_in[0], chanx_right_in[55], chanx_right_in[110], chanx_right_in[165]}),
		.sram(mux_2level_tapbuf_size6_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_23_sram_inv[0:5]),
		.out(chany_top_out[216]));

	mux_2level_tapbuf_size6 mux_bottom_track_17 (
		.in({chanx_right_in[51], chanx_right_in[106], chanx_right_in[161], chanx_right_in[216], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size6_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_24_sram_inv[0:5]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size6 mux_bottom_track_25 (
		.in({chanx_right_in[50], chanx_right_in[105], chanx_right_in[160], chanx_right_in[215], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size6_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_25_sram_inv[0:5]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size6 mux_bottom_track_33 (
		.in({chanx_right_in[49], chanx_right_in[104], chanx_right_in[159], chanx_right_in[214], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size6_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_26_sram_inv[0:5]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size6 mux_bottom_track_41 (
		.in({chanx_right_in[48], chanx_right_in[103], chanx_right_in[158], chanx_right_in[213], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size6_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_27_sram_inv[0:5]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size6 mux_bottom_track_49 (
		.in({chanx_right_in[47], chanx_right_in[102], chanx_right_in[157], chanx_right_in[212], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size6_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size6_28_sram_inv[0:5]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size6_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_0_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_1_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_2_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_3_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_4_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_5_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_6_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_7_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_8_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_9_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_10_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_11_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_12_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_13_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_14_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_15_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_16_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_17_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_18_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_19_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_20_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_376 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_21_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_22_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_top_track_432 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_23_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_24_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_25_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_26_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_27_sram_inv[0:5]));

	mux_2level_tapbuf_size6_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size6_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size6_28_sram_inv[0:5]));

	mux_2level_tapbuf_size5 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[14], chanx_right_in[69], chanx_right_in[124], chanx_right_in[179]}),
		.sram(mux_2level_tapbuf_size5_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_0_sram_inv[0:5]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size5 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[15], chanx_right_in[70], chanx_right_in[125], chanx_right_in[180]}),
		.sram(mux_2level_tapbuf_size5_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_1_sram_inv[0:5]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size5 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[16], chanx_right_in[71], chanx_right_in[126], chanx_right_in[181]}),
		.sram(mux_2level_tapbuf_size5_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_2_sram_inv[0:5]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size5 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[17], chanx_right_in[72], chanx_right_in[127], chanx_right_in[182]}),
		.sram(mux_2level_tapbuf_size5_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_3_sram_inv[0:5]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size5 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[18], chanx_right_in[73], chanx_right_in[128], chanx_right_in[183]}),
		.sram(mux_2level_tapbuf_size5_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_4_sram_inv[0:5]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size5 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[23], chanx_right_in[78], chanx_right_in[133], chanx_right_in[188]}),
		.sram(mux_2level_tapbuf_size5_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_5_sram_inv[0:5]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size5 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[24], chanx_right_in[79], chanx_right_in[134], chanx_right_in[189]}),
		.sram(mux_2level_tapbuf_size5_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_6_sram_inv[0:5]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size5 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[25], chanx_right_in[80], chanx_right_in[135], chanx_right_in[190]}),
		.sram(mux_2level_tapbuf_size5_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_7_sram_inv[0:5]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size5 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[26], chanx_right_in[81], chanx_right_in[136], chanx_right_in[191]}),
		.sram(mux_2level_tapbuf_size5_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_8_sram_inv[0:5]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size5 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[27], chanx_right_in[82], chanx_right_in[137], chanx_right_in[192]}),
		.sram(mux_2level_tapbuf_size5_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_9_sram_inv[0:5]),
		.out(chany_top_out[104]));

	mux_2level_tapbuf_size5 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[32], chanx_right_in[87], chanx_right_in[142], chanx_right_in[197]}),
		.sram(mux_2level_tapbuf_size5_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_10_sram_inv[0:5]),
		.out(chany_top_out[124]));

	mux_2level_tapbuf_size5 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[33], chanx_right_in[88], chanx_right_in[143], chanx_right_in[198]}),
		.sram(mux_2level_tapbuf_size5_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_11_sram_inv[0:5]),
		.out(chany_top_out[128]));

	mux_2level_tapbuf_size5 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[34], chanx_right_in[89], chanx_right_in[144], chanx_right_in[199]}),
		.sram(mux_2level_tapbuf_size5_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_12_sram_inv[0:5]),
		.out(chany_top_out[132]));

	mux_2level_tapbuf_size5 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[35], chanx_right_in[90], chanx_right_in[145], chanx_right_in[200]}),
		.sram(mux_2level_tapbuf_size5_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_13_sram_inv[0:5]),
		.out(chany_top_out[136]));

	mux_2level_tapbuf_size5 mux_top_track_280 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[36], chanx_right_in[91], chanx_right_in[146], chanx_right_in[201]}),
		.sram(mux_2level_tapbuf_size5_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_14_sram_inv[0:5]),
		.out(chany_top_out[140]));

	mux_2level_tapbuf_size5 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[41], chanx_right_in[96], chanx_right_in[151], chanx_right_in[206]}),
		.sram(mux_2level_tapbuf_size5_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_15_sram_inv[0:5]),
		.out(chany_top_out[160]));

	mux_2level_tapbuf_size5 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[42], chanx_right_in[97], chanx_right_in[152], chanx_right_in[207]}),
		.sram(mux_2level_tapbuf_size5_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_16_sram_inv[0:5]),
		.out(chany_top_out[164]));

	mux_2level_tapbuf_size5 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[43], chanx_right_in[98], chanx_right_in[153], chanx_right_in[208]}),
		.sram(mux_2level_tapbuf_size5_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_17_sram_inv[0:5]),
		.out(chany_top_out[168]));

	mux_2level_tapbuf_size5 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[44], chanx_right_in[99], chanx_right_in[154], chanx_right_in[209]}),
		.sram(mux_2level_tapbuf_size5_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_18_sram_inv[0:5]),
		.out(chany_top_out[172]));

	mux_2level_tapbuf_size5 mux_top_track_352 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[45], chanx_right_in[100], chanx_right_in[155], chanx_right_in[210]}),
		.sram(mux_2level_tapbuf_size5_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_19_sram_inv[0:5]),
		.out(chany_top_out[176]));

	mux_2level_tapbuf_size5 mux_top_track_392 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[50], chanx_right_in[105], chanx_right_in[160], chanx_right_in[215]}),
		.sram(mux_2level_tapbuf_size5_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_20_sram_inv[0:5]),
		.out(chany_top_out[196]));

	mux_2level_tapbuf_size5 mux_top_track_400 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[51], chanx_right_in[106], chanx_right_in[161], chanx_right_in[216]}),
		.sram(mux_2level_tapbuf_size5_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_21_sram_inv[0:5]),
		.out(chany_top_out[200]));

	mux_2level_tapbuf_size5 mux_right_track_108 (
		.in({chany_top_in[70], chany_top_in[215], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[214]}),
		.sram(mux_2level_tapbuf_size5_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_22_sram_inv[0:5]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size5 mux_bottom_track_1 (
		.in({chanx_right_in[53], chanx_right_in[108], chanx_right_in[163], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_23_sram_inv[0:5]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size5 mux_bottom_track_9 (
		.in({chanx_right_in[52], chanx_right_in[107], chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_24_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_24_sram_inv[0:5]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size5 mux_bottom_track_57 (
		.in({chanx_right_in[46], chanx_right_in[101], chanx_right_in[156], chanx_right_in[211], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_25_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_25_sram_inv[0:5]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size5 mux_bottom_track_73 (
		.in({chanx_right_in[44], chanx_right_in[99], chanx_right_in[154], chanx_right_in[209], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_26_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_26_sram_inv[0:5]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size5 mux_bottom_track_81 (
		.in({chanx_right_in[43], chanx_right_in[98], chanx_right_in[153], chanx_right_in[208], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_27_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_27_sram_inv[0:5]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size5 mux_bottom_track_89 (
		.in({chanx_right_in[42], chanx_right_in[97], chanx_right_in[152], chanx_right_in[207], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_28_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_28_sram_inv[0:5]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size5 mux_bottom_track_97 (
		.in({chanx_right_in[41], chanx_right_in[96], chanx_right_in[151], chanx_right_in[206], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_29_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_29_sram_inv[0:5]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size5 mux_bottom_track_105 (
		.in({chanx_right_in[40], chanx_right_in[95], chanx_right_in[150], chanx_right_in[205], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_30_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_30_sram_inv[0:5]),
		.out(chany_bottom_out[52]));

	mux_2level_tapbuf_size5 mux_bottom_track_113 (
		.in({chanx_right_in[39], chanx_right_in[94], chanx_right_in[149], chanx_right_in[204], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_31_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_31_sram_inv[0:5]),
		.out(chany_bottom_out[56]));

	mux_2level_tapbuf_size5 mux_bottom_track_121 (
		.in({chanx_right_in[38], chanx_right_in[93], chanx_right_in[148], chanx_right_in[203], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_32_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_32_sram_inv[0:5]),
		.out(chany_bottom_out[60]));

	mux_2level_tapbuf_size5 mux_bottom_track_129 (
		.in({chanx_right_in[37], chanx_right_in[92], chanx_right_in[147], chanx_right_in[202], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_33_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_33_sram_inv[0:5]),
		.out(chany_bottom_out[64]));

	mux_2level_tapbuf_size5 mux_bottom_track_145 (
		.in({chanx_right_in[35], chanx_right_in[90], chanx_right_in[145], chanx_right_in[200], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_34_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_34_sram_inv[0:5]),
		.out(chany_bottom_out[72]));

	mux_2level_tapbuf_size5 mux_bottom_track_153 (
		.in({chanx_right_in[34], chanx_right_in[89], chanx_right_in[144], chanx_right_in[199], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_35_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_35_sram_inv[0:5]),
		.out(chany_bottom_out[76]));

	mux_2level_tapbuf_size5 mux_bottom_track_161 (
		.in({chanx_right_in[33], chanx_right_in[88], chanx_right_in[143], chanx_right_in[198], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_36_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_36_sram_inv[0:5]),
		.out(chany_bottom_out[80]));

	mux_2level_tapbuf_size5 mux_bottom_track_169 (
		.in({chanx_right_in[32], chanx_right_in[87], chanx_right_in[142], chanx_right_in[197], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_37_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_37_sram_inv[0:5]),
		.out(chany_bottom_out[84]));

	mux_2level_tapbuf_size5 mux_bottom_track_177 (
		.in({chanx_right_in[31], chanx_right_in[86], chanx_right_in[141], chanx_right_in[196], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_38_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_38_sram_inv[0:5]),
		.out(chany_bottom_out[88]));

	mux_2level_tapbuf_size5 mux_bottom_track_185 (
		.in({chanx_right_in[30], chanx_right_in[85], chanx_right_in[140], chanx_right_in[195], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_39_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_39_sram_inv[0:5]),
		.out(chany_bottom_out[92]));

	mux_2level_tapbuf_size5 mux_bottom_track_193 (
		.in({chanx_right_in[29], chanx_right_in[84], chanx_right_in[139], chanx_right_in[194], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_40_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_40_sram_inv[0:5]),
		.out(chany_bottom_out[96]));

	mux_2level_tapbuf_size5 mux_bottom_track_201 (
		.in({chanx_right_in[28], chanx_right_in[83], chanx_right_in[138], chanx_right_in[193], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_41_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_41_sram_inv[0:5]),
		.out(chany_bottom_out[100]));

	mux_2level_tapbuf_size5 mux_bottom_track_217 (
		.in({chanx_right_in[26], chanx_right_in[81], chanx_right_in[136], chanx_right_in[191], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_42_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_42_sram_inv[0:5]),
		.out(chany_bottom_out[108]));

	mux_2level_tapbuf_size5 mux_bottom_track_225 (
		.in({chanx_right_in[25], chanx_right_in[80], chanx_right_in[135], chanx_right_in[190], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_43_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_43_sram_inv[0:5]),
		.out(chany_bottom_out[112]));

	mux_2level_tapbuf_size5 mux_bottom_track_233 (
		.in({chanx_right_in[24], chanx_right_in[79], chanx_right_in[134], chanx_right_in[189], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_44_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_44_sram_inv[0:5]),
		.out(chany_bottom_out[116]));

	mux_2level_tapbuf_size5 mux_bottom_track_241 (
		.in({chanx_right_in[23], chanx_right_in[78], chanx_right_in[133], chanx_right_in[188], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_45_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_45_sram_inv[0:5]),
		.out(chany_bottom_out[120]));

	mux_2level_tapbuf_size5 mux_bottom_track_249 (
		.in({chanx_right_in[22], chanx_right_in[77], chanx_right_in[132], chanx_right_in[187], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_46_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_46_sram_inv[0:5]),
		.out(chany_bottom_out[124]));

	mux_2level_tapbuf_size5 mux_bottom_track_257 (
		.in({chanx_right_in[21], chanx_right_in[76], chanx_right_in[131], chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_47_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_47_sram_inv[0:5]),
		.out(chany_bottom_out[128]));

	mux_2level_tapbuf_size5 mux_bottom_track_265 (
		.in({chanx_right_in[20], chanx_right_in[75], chanx_right_in[130], chanx_right_in[185], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_48_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_48_sram_inv[0:5]),
		.out(chany_bottom_out[132]));

	mux_2level_tapbuf_size5 mux_bottom_track_273 (
		.in({chanx_right_in[19], chanx_right_in[74], chanx_right_in[129], chanx_right_in[184], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_49_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_49_sram_inv[0:5]),
		.out(chany_bottom_out[136]));

	mux_2level_tapbuf_size5 mux_bottom_track_289 (
		.in({chanx_right_in[17], chanx_right_in[72], chanx_right_in[127], chanx_right_in[182], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_50_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_50_sram_inv[0:5]),
		.out(chany_bottom_out[144]));

	mux_2level_tapbuf_size5 mux_bottom_track_297 (
		.in({chanx_right_in[16], chanx_right_in[71], chanx_right_in[126], chanx_right_in[181], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_51_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_51_sram_inv[0:5]),
		.out(chany_bottom_out[148]));

	mux_2level_tapbuf_size5 mux_bottom_track_305 (
		.in({chanx_right_in[15], chanx_right_in[70], chanx_right_in[125], chanx_right_in[180], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_52_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_52_sram_inv[0:5]),
		.out(chany_bottom_out[152]));

	mux_2level_tapbuf_size5 mux_bottom_track_313 (
		.in({chanx_right_in[14], chanx_right_in[69], chanx_right_in[124], chanx_right_in[179], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_53_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_53_sram_inv[0:5]),
		.out(chany_bottom_out[156]));

	mux_2level_tapbuf_size5 mux_bottom_track_321 (
		.in({chanx_right_in[13], chanx_right_in[68], chanx_right_in[123], chanx_right_in[178], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_54_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_54_sram_inv[0:5]),
		.out(chany_bottom_out[160]));

	mux_2level_tapbuf_size5 mux_bottom_track_329 (
		.in({chanx_right_in[12], chanx_right_in[67], chanx_right_in[122], chanx_right_in[177], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_55_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_55_sram_inv[0:5]),
		.out(chany_bottom_out[164]));

	mux_2level_tapbuf_size5 mux_bottom_track_337 (
		.in({chanx_right_in[11], chanx_right_in[66], chanx_right_in[121], chanx_right_in[176], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_56_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_56_sram_inv[0:5]),
		.out(chany_bottom_out[168]));

	mux_2level_tapbuf_size5 mux_bottom_track_345 (
		.in({chanx_right_in[10], chanx_right_in[65], chanx_right_in[120], chanx_right_in[175], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_57_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_57_sram_inv[0:5]),
		.out(chany_bottom_out[172]));

	mux_2level_tapbuf_size5 mux_bottom_track_361 (
		.in({chanx_right_in[8], chanx_right_in[63], chanx_right_in[118], chanx_right_in[173], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_58_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_58_sram_inv[0:5]),
		.out(chany_bottom_out[180]));

	mux_2level_tapbuf_size5 mux_bottom_track_369 (
		.in({chanx_right_in[7], chanx_right_in[62], chanx_right_in[117], chanx_right_in[172], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_59_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_59_sram_inv[0:5]),
		.out(chany_bottom_out[184]));

	mux_2level_tapbuf_size5 mux_bottom_track_377 (
		.in({chanx_right_in[6], chanx_right_in[61], chanx_right_in[116], chanx_right_in[171], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_60_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_60_sram_inv[0:5]),
		.out(chany_bottom_out[188]));

	mux_2level_tapbuf_size5 mux_bottom_track_385 (
		.in({chanx_right_in[5], chanx_right_in[60], chanx_right_in[115], chanx_right_in[170], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_61_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_61_sram_inv[0:5]),
		.out(chany_bottom_out[192]));

	mux_2level_tapbuf_size5 mux_bottom_track_393 (
		.in({chanx_right_in[4], chanx_right_in[59], chanx_right_in[114], chanx_right_in[169], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_62_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_62_sram_inv[0:5]),
		.out(chany_bottom_out[196]));

	mux_2level_tapbuf_size5 mux_bottom_track_401 (
		.in({chanx_right_in[3], chanx_right_in[58], chanx_right_in[113], chanx_right_in[168], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_63_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_63_sram_inv[0:5]),
		.out(chany_bottom_out[200]));

	mux_2level_tapbuf_size5 mux_bottom_track_409 (
		.in({chanx_right_in[2], chanx_right_in[57], chanx_right_in[112], chanx_right_in[167], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_64_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_64_sram_inv[0:5]),
		.out(chany_bottom_out[204]));

	mux_2level_tapbuf_size5 mux_bottom_track_417 (
		.in({chanx_right_in[1], chanx_right_in[56], chanx_right_in[111], chanx_right_in[166], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size5_65_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size5_65_sram_inv[0:5]),
		.out(chany_bottom_out[208]));

	mux_2level_tapbuf_size5_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_0_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_1_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_2_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_3_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_4_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_5_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_6_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_7_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_8_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_9_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_10_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_11_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_12_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_13_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_14_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_15_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_16_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_17_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_18_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_19_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_20_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_top_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_21_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_22_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_23_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_24_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_24_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_25_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_25_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_26_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_26_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_27_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_27_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_28_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_28_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_29_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_29_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_105 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_30_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_30_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_113 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_31_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_31_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_121 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_32_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_32_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_129 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_33_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_33_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_145 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_34_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_34_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_153 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_35_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_35_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_161 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_36_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_36_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_169 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_37_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_37_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_177 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_38_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_38_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_185 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_39_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_39_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_193 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_40_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_40_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_201 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_41_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_41_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_217 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_42_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_42_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_225 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_43_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_43_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_233 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_44_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_44_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_241 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_45_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_45_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_249 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_46_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_46_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_257 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_47_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_47_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_265 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_48_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_48_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_273 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_49_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_49_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_289 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_50_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_50_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_297 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_51_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_51_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_305 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_52_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_52_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_313 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_53_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_53_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_321 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_54_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_54_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_329 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_55_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_55_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_337 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_56_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_56_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_345 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_57_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_57_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_361 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_58_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_58_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_369 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_59_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_59_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_377 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_60_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_60_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_385 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_61_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_61_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_393 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_62_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_62_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_401 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_63_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_63_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_409 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_64_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_64_sram_inv[0:5]));

	mux_2level_tapbuf_size5_mem mem_bottom_track_417 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size5_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size5_65_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size5_65_sram_inv[0:5]));

	mux_2level_tapbuf_size4 mux_top_track_408 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[52], chanx_right_in[107], chanx_right_in[162]}),
		.sram(mux_2level_tapbuf_size4_0_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_0_sram_inv[0:5]),
		.out(chany_top_out[204]));

	mux_2level_tapbuf_size4 mux_top_track_416 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[53], chanx_right_in[108], chanx_right_in[163]}),
		.sram(mux_2level_tapbuf_size4_1_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_1_sram_inv[0:5]),
		.out(chany_top_out[208]));

	mux_2level_tapbuf_size4 mux_top_track_424 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[54], chanx_right_in[109], chanx_right_in[164]}),
		.sram(mux_2level_tapbuf_size4_2_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_2_sram_inv[0:5]),
		.out(chany_top_out[212]));

	mux_2level_tapbuf_size4 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size4_3_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_3_sram_inv[0:5]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size4 mux_right_track_110 (
		.in({chany_top_in[72], chany_top_in[216], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[213]}),
		.sram(mux_2level_tapbuf_size4_4_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_4_sram_inv[0:5]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size4 mux_right_track_126 (
		.in({chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[202]}),
		.sram(mux_2level_tapbuf_size4_5_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_5_sram_inv[0:5]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size4 mux_right_track_128 (
		.in({chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[201]}),
		.sram(mux_2level_tapbuf_size4_6_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_6_sram_inv[0:5]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size4 mux_right_track_146 (
		.in({chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[189]}),
		.sram(mux_2level_tapbuf_size4_7_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_7_sram_inv[0:5]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size4 mux_right_track_148 (
		.in({chany_top_in[97], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[188]}),
		.sram(mux_2level_tapbuf_size4_8_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_8_sram_inv[0:5]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size4 mux_right_track_166 (
		.in({chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[176]}),
		.sram(mux_2level_tapbuf_size4_9_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_9_sram_inv[0:5]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size4 mux_right_track_288 (
		.in({chany_top_in[190], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[94]}),
		.sram(mux_2level_tapbuf_size4_10_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_10_sram_inv[0:5]),
		.out(chanx_right_out[144]));

	mux_2level_tapbuf_size4 mux_right_track_306 (
		.in({chany_top_in[202], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[82]}),
		.sram(mux_2level_tapbuf_size4_11_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_11_sram_inv[0:5]),
		.out(chanx_right_out[153]));

	mux_2level_tapbuf_size4 mux_right_track_308 (
		.in({chany_top_in[204], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[81]}),
		.sram(mux_2level_tapbuf_size4_12_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_12_sram_inv[0:5]),
		.out(chanx_right_out[154]));

	mux_2level_tapbuf_size4 mux_right_track_324 (
		.in({chany_top_in[214], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[70], chany_bottom_in[215]}),
		.sram(mux_2level_tapbuf_size4_13_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_13_sram_inv[0:5]),
		.out(chanx_right_out[162]));

	mux_2level_tapbuf_size4 mux_right_track_326 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[69], chany_bottom_in[211]}),
		.sram(mux_2level_tapbuf_size4_14_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_14_sram_inv[0:5]),
		.out(chanx_right_out[163]));

	mux_2level_tapbuf_size4 mux_right_track_328 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[68], chany_bottom_in[207]}),
		.sram(mux_2level_tapbuf_size4_15_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_15_sram_inv[0:5]),
		.out(chanx_right_out[164]));

	mux_2level_tapbuf_size4 mux_right_track_346 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[56], chany_bottom_in[171]}),
		.sram(mux_2level_tapbuf_size4_16_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_16_sram_inv[0:5]),
		.out(chanx_right_out[173]));

	mux_2level_tapbuf_size4 mux_bottom_track_65 (
		.in({chanx_right_in[45], chanx_right_in[100], chanx_right_in[155], chanx_right_in[210]}),
		.sram(mux_2level_tapbuf_size4_17_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_17_sram_inv[0:5]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size4 mux_bottom_track_137 (
		.in({chanx_right_in[36], chanx_right_in[91], chanx_right_in[146], chanx_right_in[201]}),
		.sram(mux_2level_tapbuf_size4_18_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_18_sram_inv[0:5]),
		.out(chany_bottom_out[68]));

	mux_2level_tapbuf_size4 mux_bottom_track_209 (
		.in({chanx_right_in[27], chanx_right_in[82], chanx_right_in[137], chanx_right_in[192]}),
		.sram(mux_2level_tapbuf_size4_19_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_19_sram_inv[0:5]),
		.out(chany_bottom_out[104]));

	mux_2level_tapbuf_size4 mux_bottom_track_281 (
		.in({chanx_right_in[18], chanx_right_in[73], chanx_right_in[128], chanx_right_in[183]}),
		.sram(mux_2level_tapbuf_size4_20_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_20_sram_inv[0:5]),
		.out(chany_bottom_out[140]));

	mux_2level_tapbuf_size4 mux_bottom_track_353 (
		.in({chanx_right_in[9], chanx_right_in[64], chanx_right_in[119], chanx_right_in[174]}),
		.sram(mux_2level_tapbuf_size4_21_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_21_sram_inv[0:5]),
		.out(chany_bottom_out[176]));

	mux_2level_tapbuf_size4 mux_bottom_track_425 (
		.in({chanx_right_in[0], chanx_right_in[55], chanx_right_in[110], chanx_right_in[165]}),
		.sram(mux_2level_tapbuf_size4_22_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_22_sram_inv[0:5]),
		.out(chany_bottom_out[212]));

	mux_2level_tapbuf_size4 mux_bottom_track_433 (
		.in({chanx_right_in[54], chanx_right_in[109], chanx_right_in[164], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size4_23_sram[0:5]),
		.sram_inv(mux_2level_tapbuf_size4_23_sram_inv[0:5]),
		.out(chany_bottom_out[216]));

	mux_2level_tapbuf_size4_mem mem_top_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_0_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_0_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_top_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_1_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_1_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_top_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_2_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_2_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_3_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_3_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_4_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_4_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_5_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_5_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_6_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_6_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_7_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_7_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_8_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_8_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_9_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_9_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_288 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_10_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_10_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_306 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_11_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_11_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_12_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_12_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_324 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_13_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_13_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_326 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_14_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_14_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_328 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_15_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_15_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_right_track_346 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_16_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_16_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_17_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_17_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_137 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_18_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_18_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_209 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_19_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_19_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_281 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_20_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_20_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_353 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_21_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_21_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_425 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size5_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size4_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_22_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_22_sram_inv[0:5]));

	mux_2level_tapbuf_size4_mem mem_bottom_track_433 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_22_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size4_23_sram[0:5]),
		.mem_outb(mux_2level_tapbuf_size4_23_sram_inv[0:5]));

	mux_2level_tapbuf_size2 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size2 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size2 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size2 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size2 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size2 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size2 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size2 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size2 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size2 mux_right_track_42 (
		.in({chany_top_in[26], chany_top_in[83]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size2 mux_right_track_44 (
		.in({chany_top_in[28], chany_top_in[87]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size2 mux_right_track_50 (
		.in({chany_top_in[32], chany_top_in[99]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size2 mux_right_track_52 (
		.in({chany_top_in[33], chany_top_in[103]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size2 mux_right_track_60 (
		.in({chany_top_in[38], chany_top_in[119]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size2 mux_right_track_62 (
		.in({chany_top_in[40], chany_top_in[123]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size2 mux_right_track_64 (
		.in({chany_top_in[41], chany_top_in[127]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size2 mux_right_track_70 (
		.in({chany_top_in[45], chany_top_in[139]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_2level_tapbuf_size2 mux_right_track_78 (
		.in({chany_top_in[50], chany_top_in[155]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size2 mux_right_track_80 (
		.in({chany_top_in[52], chany_top_in[159]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size2 mux_right_track_82 (
		.in({chany_top_in[53], chany_top_in[163]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size2 mux_right_track_84 (
		.in({chany_top_in[54], chany_top_in[167]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size2 mux_right_track_96 (
		.in({chany_top_in[62], chany_top_in[191]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size2 mux_right_track_98 (
		.in({chany_top_in[64], chany_top_in[195]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size2 mux_right_track_100 (
		.in({chany_top_in[65], chany_top_in[199]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size2 mux_right_track_102 (
		.in({chany_top_in[66], chany_top_in[203]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size2 mux_right_track_104 (
		.in({chany_top_in[68], chany_top_in[207]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size2 mux_right_track_114 (
		.in({chany_top_in[74], chany_bottom_in[210]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size2 mux_right_track_116 (
		.in({chany_top_in[76], chany_bottom_in[209]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size2 mux_right_track_118 (
		.in({chany_top_in[77], chany_bottom_in[208]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_2level_tapbuf_size2 mux_right_track_120 (
		.in({chany_top_in[78], chany_bottom_in[206]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size2 mux_right_track_122 (
		.in({chany_top_in[80], chany_bottom_in[205]}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size2 mux_right_track_124 (
		.in({chany_top_in[81], chany_bottom_in[204]}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_2level_tapbuf_size2 mux_right_track_132 (
		.in({chany_top_in[86], chany_bottom_in[198]}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size2 mux_right_track_134 (
		.in({chany_top_in[88], chany_bottom_in[197]}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size2 mux_right_track_136 (
		.in({chany_top_in[89], chany_bottom_in[196]}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size2 mux_right_track_138 (
		.in({chany_top_in[90], chany_bottom_in[194]}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size2 mux_right_track_140 (
		.in({chany_top_in[92], chany_bottom_in[193]}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size2 mux_right_track_142 (
		.in({chany_top_in[93], chany_bottom_in[192]}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_2level_tapbuf_size2 mux_right_track_150 (
		.in({chany_top_in[98], chany_bottom_in[186]}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size2 mux_right_track_152 (
		.in({chany_top_in[100], chany_bottom_in[185]}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size2 mux_right_track_154 (
		.in({chany_top_in[101], chany_bottom_in[184]}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size2 mux_right_track_156 (
		.in({chany_top_in[102], chany_bottom_in[182]}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size2 mux_right_track_158 (
		.in({chany_top_in[104], chany_bottom_in[181]}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_2level_tapbuf_size2 mux_right_track_160 (
		.in({chany_top_in[105], chany_bottom_in[180]}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_2level_tapbuf_size2 mux_right_track_170 (
		.in({chany_top_in[112], chany_bottom_in[173]}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size2 mux_right_track_172 (
		.in({chany_top_in[113], chany_bottom_in[172]}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size2 mux_right_track_174 (
		.in({chany_top_in[114], chany_bottom_in[170]}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size2 mux_right_track_176 (
		.in({chany_top_in[116], chany_bottom_in[169]}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size2 mux_right_track_178 (
		.in({chany_top_in[117], chany_bottom_in[168]}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_2level_tapbuf_size2 mux_right_track_190 (
		.in({chany_top_in[125], chany_bottom_in[160]}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size2 mux_right_track_192 (
		.in({chany_top_in[126], chany_bottom_in[158]}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size2 mux_right_track_194 (
		.in({chany_top_in[128], chany_bottom_in[157]}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size2 mux_right_track_196 (
		.in({chany_top_in[129], chany_bottom_in[156]}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_2level_tapbuf_size2 mux_right_track_204 (
		.in({chany_top_in[134], chany_bottom_in[150]}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size2 mux_right_track_210 (
		.in({chany_top_in[138], chany_bottom_in[146]}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_2level_tapbuf_size2 mux_right_track_212 (
		.in({chany_top_in[140], chany_bottom_in[145]}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size2 mux_right_track_214 (
		.in({chany_top_in[141], chany_bottom_in[144]}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_2level_tapbuf_size2 mux_right_track_222 (
		.in({chany_top_in[146], chany_bottom_in[138]}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_2level_tapbuf_size2 mux_right_track_224 (
		.in({chany_top_in[148], chany_bottom_in[137]}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_2level_tapbuf_size2 mux_right_track_230 (
		.in({chany_top_in[152], chany_bottom_in[133]}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_2level_tapbuf_size2 mux_right_track_232 (
		.in({chany_top_in[153], chany_bottom_in[132]}),
		.sram(mux_2level_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_2level_tapbuf_size2 mux_right_track_240 (
		.in({chany_top_in[158], chany_bottom_in[126]}),
		.sram(mux_2level_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_2level_tapbuf_size2 mux_right_track_242 (
		.in({chany_top_in[160], chany_bottom_in[125]}),
		.sram(mux_2level_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_2level_tapbuf_size2 mux_right_track_244 (
		.in({chany_top_in[161], chany_bottom_in[124]}),
		.sram(mux_2level_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size2 mux_right_track_250 (
		.in({chany_top_in[165], chany_bottom_in[120]}),
		.sram(mux_2level_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_2level_tapbuf_size2 mux_right_track_258 (
		.in({chany_top_in[170], chany_bottom_in[114]}),
		.sram(mux_2level_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_2level_tapbuf_size2 mux_right_track_260 (
		.in({chany_top_in[172], chany_bottom_in[113]}),
		.sram(mux_2level_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size2 mux_right_track_262 (
		.in({chany_top_in[173], chany_bottom_in[112]}),
		.sram(mux_2level_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_2level_tapbuf_size2 mux_right_track_264 (
		.in({chany_top_in[174], chany_bottom_in[110]}),
		.sram(mux_2level_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_2level_tapbuf_size2 mux_right_track_276 (
		.in({chany_top_in[182], chany_bottom_in[102]}),
		.sram(mux_2level_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_2level_tapbuf_size2 mux_right_track_278 (
		.in({chany_top_in[184], chany_bottom_in[101]}),
		.sram(mux_2level_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_2level_tapbuf_size2 mux_right_track_280 (
		.in({chany_top_in[185], chany_bottom_in[100]}),
		.sram(mux_2level_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_2level_tapbuf_size2 mux_right_track_282 (
		.in({chany_top_in[186], chany_bottom_in[98]}),
		.sram(mux_2level_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_2level_tapbuf_size2 mux_right_track_284 (
		.in({chany_top_in[188], chany_bottom_in[97]}),
		.sram(mux_2level_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size2 mux_right_track_294 (
		.in({chany_top_in[194], chany_bottom_in[90]}),
		.sram(mux_2level_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_2level_tapbuf_size2 mux_right_track_296 (
		.in({chany_top_in[196], chany_bottom_in[89]}),
		.sram(mux_2level_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_2level_tapbuf_size2 mux_right_track_298 (
		.in({chany_top_in[197], chany_bottom_in[88]}),
		.sram(mux_2level_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_2level_tapbuf_size2 mux_right_track_300 (
		.in({chany_top_in[198], chany_bottom_in[86]}),
		.sram(mux_2level_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_2level_tapbuf_size2 mux_right_track_302 (
		.in({chany_top_in[200], chany_bottom_in[85]}),
		.sram(mux_2level_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_2level_tapbuf_size2 mux_right_track_304 (
		.in({chany_top_in[201], chany_bottom_in[84]}),
		.sram(mux_2level_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_right_out[152]));

	mux_2level_tapbuf_size2 mux_right_track_312 (
		.in({chany_top_in[206], chany_bottom_in[78]}),
		.sram(mux_2level_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_2level_tapbuf_size2 mux_right_track_314 (
		.in({chany_top_in[208], chany_bottom_in[77]}),
		.sram(mux_2level_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_2level_tapbuf_size2 mux_right_track_316 (
		.in({chany_top_in[209], chany_bottom_in[76]}),
		.sram(mux_2level_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_2level_tapbuf_size2 mux_right_track_318 (
		.in({chany_top_in[210], chany_bottom_in[74]}),
		.sram(mux_2level_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_83_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_2level_tapbuf_size2 mux_right_track_320 (
		.in({chany_top_in[212], chany_bottom_in[73]}),
		.sram(mux_2level_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_84_sram_inv[0:1]),
		.out(chanx_right_out[160]));

	mux_2level_tapbuf_size2 mux_right_track_330 (
		.in({chany_bottom_in[66], chany_bottom_in[203]}),
		.sram(mux_2level_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_85_sram_inv[0:1]),
		.out(chanx_right_out[165]));

	mux_2level_tapbuf_size2 mux_right_track_332 (
		.in({chany_bottom_in[65], chany_bottom_in[199]}),
		.sram(mux_2level_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_86_sram_inv[0:1]),
		.out(chanx_right_out[166]));

	mux_2level_tapbuf_size2 mux_right_track_334 (
		.in({chany_bottom_in[64], chany_bottom_in[195]}),
		.sram(mux_2level_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_87_sram_inv[0:1]),
		.out(chanx_right_out[167]));

	mux_2level_tapbuf_size2 mux_right_track_336 (
		.in({chany_bottom_in[62], chany_bottom_in[191]}),
		.sram(mux_2level_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_88_sram_inv[0:1]),
		.out(chanx_right_out[168]));

	mux_2level_tapbuf_size2 mux_right_track_338 (
		.in({chany_bottom_in[61], chany_bottom_in[187]}),
		.sram(mux_2level_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_89_sram_inv[0:1]),
		.out(chanx_right_out[169]));

	mux_2level_tapbuf_size2 mux_right_track_340 (
		.in({chany_bottom_in[60], chany_bottom_in[183]}),
		.sram(mux_2level_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_90_sram_inv[0:1]),
		.out(chanx_right_out[170]));

	mux_2level_tapbuf_size2 mux_right_track_350 (
		.in({chany_bottom_in[53], chany_bottom_in[163]}),
		.sram(mux_2level_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_91_sram_inv[0:1]),
		.out(chanx_right_out[175]));

	mux_2level_tapbuf_size2 mux_right_track_352 (
		.in({chany_bottom_in[52], chany_bottom_in[159]}),
		.sram(mux_2level_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_92_sram_inv[0:1]),
		.out(chanx_right_out[176]));

	mux_2level_tapbuf_size2 mux_right_track_354 (
		.in({chany_bottom_in[50], chany_bottom_in[155]}),
		.sram(mux_2level_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_93_sram_inv[0:1]),
		.out(chanx_right_out[177]));

	mux_2level_tapbuf_size2 mux_right_track_356 (
		.in({chany_bottom_in[49], chany_bottom_in[151]}),
		.sram(mux_2level_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_94_sram_inv[0:1]),
		.out(chanx_right_out[178]));

	mux_2level_tapbuf_size2 mux_right_track_358 (
		.in({chany_bottom_in[48], chany_bottom_in[147]}),
		.sram(mux_2level_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_95_sram_inv[0:1]),
		.out(chanx_right_out[179]));

	mux_2level_tapbuf_size2 mux_right_track_370 (
		.in({chany_bottom_in[40], chany_bottom_in[123]}),
		.sram(mux_2level_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_96_sram_inv[0:1]),
		.out(chanx_right_out[185]));

	mux_2level_tapbuf_size2 mux_right_track_372 (
		.in({chany_bottom_in[38], chany_bottom_in[119]}),
		.sram(mux_2level_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_97_sram_inv[0:1]),
		.out(chanx_right_out[186]));

	mux_2level_tapbuf_size2 mux_right_track_374 (
		.in({chany_bottom_in[37], chany_bottom_in[115]}),
		.sram(mux_2level_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_98_sram_inv[0:1]),
		.out(chanx_right_out[187]));

	mux_2level_tapbuf_size2 mux_right_track_376 (
		.in({chany_bottom_in[36], chany_bottom_in[111]}),
		.sram(mux_2level_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_99_sram_inv[0:1]),
		.out(chanx_right_out[188]));

	mux_2level_tapbuf_size2 mux_right_track_384 (
		.in({chany_bottom_in[30], chany_bottom_in[95]}),
		.sram(mux_2level_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_100_sram_inv[0:1]),
		.out(chanx_right_out[192]));

	mux_2level_tapbuf_size2 mux_right_track_390 (
		.in({chany_bottom_in[26], chany_bottom_in[83]}),
		.sram(mux_2level_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_101_sram_inv[0:1]),
		.out(chanx_right_out[195]));

	mux_2level_tapbuf_size2 mux_right_track_392 (
		.in({chany_bottom_in[25], chany_bottom_in[79]}),
		.sram(mux_2level_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_102_sram_inv[0:1]),
		.out(chanx_right_out[196]));

	mux_2level_tapbuf_size2 mux_right_track_394 (
		.in({chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_2level_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_103_sram_inv[0:1]),
		.out(chanx_right_out[197]));

	mux_2level_tapbuf_size2 mux_right_track_402 (
		.in({chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_2level_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_104_sram_inv[0:1]),
		.out(chanx_right_out[201]));

	mux_2level_tapbuf_size2 mux_right_track_404 (
		.in({chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_2level_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_105_sram_inv[0:1]),
		.out(chanx_right_out[202]));

	mux_2level_tapbuf_size2 mux_right_track_410 (
		.in({chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_2level_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_106_sram_inv[0:1]),
		.out(chanx_right_out[205]));

	mux_2level_tapbuf_size2 mux_right_track_412 (
		.in({chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_2level_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_107_sram_inv[0:1]),
		.out(chanx_right_out[206]));

	mux_2level_tapbuf_size2 mux_right_track_420 (
		.in({chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_2level_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_108_sram_inv[0:1]),
		.out(chanx_right_out[210]));

	mux_2level_tapbuf_size2 mux_right_track_422 (
		.in({chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_2level_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_109_sram_inv[0:1]),
		.out(chanx_right_out[211]));

	mux_2level_tapbuf_size2 mux_right_track_424 (
		.in({chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_2level_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_110_sram_inv[0:1]),
		.out(chanx_right_out[212]));

	mux_2level_tapbuf_size2 mux_right_track_430 (
		.in({chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_2level_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_111_sram_inv[0:1]),
		.out(chanx_right_out[215]));

	mux_2level_tapbuf_size2_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_142 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_160 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_178 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_210 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_214 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_222 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_224 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_230 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_232 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_60_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_240 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_61_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_242 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_62_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_63_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_250 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_64_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_258 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_65_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_66_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_262 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_67_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_264 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_68_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_69_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_278 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_70_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_280 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_71_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_282 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_72_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_73_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_294 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_74_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_296 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_75_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_298 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_76_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_77_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_302 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_78_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_304 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_79_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_312 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_80_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_314 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_81_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_82_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_318 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_83_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_320 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_84_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_330 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_85_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_332 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_86_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_334 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_87_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_336 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_88_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_338 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_89_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_340 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_90_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_350 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_91_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_352 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_92_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_354 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_93_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_356 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_94_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_358 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_95_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_370 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_96_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_372 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_97_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_374 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_98_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_376 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_99_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_384 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_100_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_390 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_101_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_392 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_102_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_394 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_103_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_402 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_104_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_404 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_105_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_410 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_106_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_412 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_107_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_420 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_108_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_422 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_109_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_424 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_110_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_430 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_111_sram_inv[0:1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size3 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size3 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size3 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size3 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size3 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size3 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size3 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_2level_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size3 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size3 mux_right_track_40 (
		.in({chany_top_in[25], chany_top_in[79], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size3 mux_right_track_46 (
		.in({chany_top_in[29], chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size3 mux_right_track_48 (
		.in({chany_top_in[30], chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size3 mux_right_track_54 (
		.in({chany_top_in[34], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_2level_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size3 mux_right_track_56 (
		.in({chany_top_in[36], chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size3 mux_right_track_58 (
		.in({chany_top_in[37], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size3 mux_right_track_66 (
		.in({chany_top_in[42], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size3 mux_right_track_68 (
		.in({chany_top_in[44], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size3 mux_right_track_72 (
		.in({chany_top_in[46], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_2level_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size3 mux_right_track_74 (
		.in({chany_top_in[48], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size3 mux_right_track_76 (
		.in({chany_top_in[49], chany_top_in[151], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size3 mux_right_track_86 (
		.in({chany_top_in[56], chany_top_in[171], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size3 mux_right_track_88 (
		.in({chany_top_in[57], chany_top_in[175], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(mux_2level_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size3 mux_right_track_90 (
		.in({chany_top_in[58], chany_top_in[179], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_2level_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size3 mux_right_track_92 (
		.in({chany_top_in[60], chany_top_in[183], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_2level_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size3 mux_right_track_94 (
		.in({chany_top_in[61], chany_top_in[187], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_}),
		.sram(mux_2level_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size3 mux_right_track_106 (
		.in({chany_top_in[69], chany_top_in[211], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(mux_2level_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_2level_tapbuf_size3 mux_right_track_112 (
		.in({chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[212]}),
		.sram(mux_2level_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size3 mux_right_track_130 (
		.in({chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[200]}),
		.sram(mux_2level_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size3 mux_right_track_144 (
		.in({chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[190]}),
		.sram(mux_2level_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size3 mux_right_track_162 (
		.in({chany_top_in[106], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[178]}),
		.sram(mux_2level_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size3 mux_right_track_164 (
		.in({chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[177]}),
		.sram(mux_2level_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size3 mux_right_track_168 (
		.in({chany_top_in[110], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[174]}),
		.sram(mux_2level_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size3 mux_right_track_180 (
		.in({chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[166]}),
		.sram(mux_2level_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size3 mux_right_track_182 (
		.in({chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[165]}),
		.sram(mux_2level_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size3 mux_right_track_184 (
		.in({chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[164]}),
		.sram(mux_2level_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size3 mux_right_track_186 (
		.in({chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[162]}),
		.sram(mux_2level_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size3 mux_right_track_188 (
		.in({chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[161]}),
		.sram(mux_2level_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size3 mux_right_track_198 (
		.in({chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[154]}),
		.sram(mux_2level_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_2level_tapbuf_size3 mux_right_track_200 (
		.in({chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[153]}),
		.sram(mux_2level_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size3 mux_right_track_202 (
		.in({chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[152]}),
		.sram(mux_2level_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size3 mux_right_track_206 (
		.in({chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[149]}),
		.sram(mux_2level_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_2level_tapbuf_size3 mux_right_track_208 (
		.in({chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[148]}),
		.sram(mux_2level_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_2level_tapbuf_size3 mux_right_track_216 (
		.in({chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[142]}),
		.sram(mux_2level_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_2level_tapbuf_size3 mux_right_track_218 (
		.in({chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[141]}),
		.sram(mux_2level_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_2level_tapbuf_size3 mux_right_track_220 (
		.in({chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[140]}),
		.sram(mux_2level_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size3 mux_right_track_226 (
		.in({chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[136]}),
		.sram(mux_2level_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_2level_tapbuf_size3 mux_right_track_228 (
		.in({chany_top_in[150], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[134]}),
		.sram(mux_2level_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size3 mux_right_track_234 (
		.in({chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[130]}),
		.sram(mux_2level_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_2level_tapbuf_size3 mux_right_track_236 (
		.in({chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[129]}),
		.sram(mux_2level_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_2level_tapbuf_size3 mux_right_track_238 (
		.in({chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[128]}),
		.sram(mux_2level_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_2level_tapbuf_size3 mux_right_track_246 (
		.in({chany_top_in[162], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[122]}),
		.sram(mux_2level_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_2level_tapbuf_size3 mux_right_track_248 (
		.in({chany_top_in[164], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[121]}),
		.sram(mux_2level_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_2level_tapbuf_size3 mux_right_track_252 (
		.in({chany_top_in[166], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[118]}),
		.sram(mux_2level_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size3 mux_right_track_254 (
		.in({chany_top_in[168], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[117]}),
		.sram(mux_2level_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_2level_tapbuf_size3 mux_right_track_256 (
		.in({chany_top_in[169], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[116]}),
		.sram(mux_2level_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_55_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_2level_tapbuf_size3 mux_right_track_266 (
		.in({chany_top_in[176], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[109]}),
		.sram(mux_2level_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_56_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_2level_tapbuf_size3 mux_right_track_268 (
		.in({chany_top_in[177], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[108]}),
		.sram(mux_2level_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_57_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_2level_tapbuf_size3 mux_right_track_270 (
		.in({chany_top_in[178], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[106]}),
		.sram(mux_2level_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_58_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_2level_tapbuf_size3 mux_right_track_272 (
		.in({chany_top_in[180], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[105]}),
		.sram(mux_2level_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_59_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_2level_tapbuf_size3 mux_right_track_274 (
		.in({chany_top_in[181], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[104]}),
		.sram(mux_2level_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_60_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_2level_tapbuf_size3 mux_right_track_286 (
		.in({chany_top_in[189], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[96]}),
		.sram(mux_2level_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_61_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_2level_tapbuf_size3 mux_right_track_290 (
		.in({chany_top_in[192], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[93]}),
		.sram(mux_2level_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_62_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_2level_tapbuf_size3 mux_right_track_292 (
		.in({chany_top_in[193], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[92]}),
		.sram(mux_2level_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_63_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size3 mux_right_track_310 (
		.in({chany_top_in[205], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[80]}),
		.sram(mux_2level_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_64_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_2level_tapbuf_size3 mux_right_track_322 (
		.in({chany_top_in[213], chany_bottom_in[72], chany_bottom_in[216]}),
		.sram(mux_2level_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_65_sram_inv[0:1]),
		.out(chanx_right_out[161]));

	mux_2level_tapbuf_size3 mux_right_track_342 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[58], chany_bottom_in[179]}),
		.sram(mux_2level_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_66_sram_inv[0:1]),
		.out(chanx_right_out[171]));

	mux_2level_tapbuf_size3 mux_right_track_344 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[57], chany_bottom_in[175]}),
		.sram(mux_2level_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_67_sram_inv[0:1]),
		.out(chanx_right_out[172]));

	mux_2level_tapbuf_size3 mux_right_track_348 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[54], chany_bottom_in[167]}),
		.sram(mux_2level_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_68_sram_inv[0:1]),
		.out(chanx_right_out[174]));

	mux_2level_tapbuf_size3 mux_right_track_360 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[46], chany_bottom_in[143]}),
		.sram(mux_2level_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_69_sram_inv[0:1]),
		.out(chanx_right_out[180]));

	mux_2level_tapbuf_size3 mux_right_track_362 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[45], chany_bottom_in[139]}),
		.sram(mux_2level_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_70_sram_inv[0:1]),
		.out(chanx_right_out[181]));

	mux_2level_tapbuf_size3 mux_right_track_364 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[44], chany_bottom_in[135]}),
		.sram(mux_2level_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_71_sram_inv[0:1]),
		.out(chanx_right_out[182]));

	mux_2level_tapbuf_size3 mux_right_track_366 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[42], chany_bottom_in[131]}),
		.sram(mux_2level_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_72_sram_inv[0:1]),
		.out(chanx_right_out[183]));

	mux_2level_tapbuf_size3 mux_right_track_368 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[41], chany_bottom_in[127]}),
		.sram(mux_2level_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_73_sram_inv[0:1]),
		.out(chanx_right_out[184]));

	mux_2level_tapbuf_size3 mux_right_track_378 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[34], chany_bottom_in[107]}),
		.sram(mux_2level_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_74_sram_inv[0:1]),
		.out(chanx_right_out[189]));

	mux_2level_tapbuf_size3 mux_right_track_380 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[33], chany_bottom_in[103]}),
		.sram(mux_2level_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_75_sram_inv[0:1]),
		.out(chanx_right_out[190]));

	mux_2level_tapbuf_size3 mux_right_track_382 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[32], chany_bottom_in[99]}),
		.sram(mux_2level_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_76_sram_inv[0:1]),
		.out(chanx_right_out[191]));

	mux_2level_tapbuf_size3 mux_right_track_386 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[29], chany_bottom_in[91]}),
		.sram(mux_2level_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_77_sram_inv[0:1]),
		.out(chanx_right_out[193]));

	mux_2level_tapbuf_size3 mux_right_track_388 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[28], chany_bottom_in[87]}),
		.sram(mux_2level_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_78_sram_inv[0:1]),
		.out(chanx_right_out[194]));

	mux_2level_tapbuf_size3 mux_right_track_396 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_2level_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_79_sram_inv[0:1]),
		.out(chanx_right_out[198]));

	mux_2level_tapbuf_size3 mux_right_track_398 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_2level_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_80_sram_inv[0:1]),
		.out(chanx_right_out[199]));

	mux_2level_tapbuf_size3 mux_right_track_400 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_2level_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_81_sram_inv[0:1]),
		.out(chanx_right_out[200]));

	mux_2level_tapbuf_size3 mux_right_track_406 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_2level_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_82_sram_inv[0:1]),
		.out(chanx_right_out[203]));

	mux_2level_tapbuf_size3 mux_right_track_408 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_2level_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_83_sram_inv[0:1]),
		.out(chanx_right_out[204]));

	mux_2level_tapbuf_size3 mux_right_track_414 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_2level_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_84_sram_inv[0:1]),
		.out(chanx_right_out[207]));

	mux_2level_tapbuf_size3 mux_right_track_416 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_2level_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_85_sram_inv[0:1]),
		.out(chanx_right_out[208]));

	mux_2level_tapbuf_size3 mux_right_track_418 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_2level_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_right_out[209]));

	mux_2level_tapbuf_size3 mux_right_track_426 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_2level_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_right_out[213]));

	mux_2level_tapbuf_size3 mux_right_track_428 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_2level_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_right_out[214]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_8_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_9_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_10_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_11_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_12_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_13_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_14_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_15_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_16_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_17_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_18_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_19_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_20_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_21_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_22_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_23_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_24_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_25_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_106 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_26_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_27_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_28_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_29_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_30_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_31_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_32_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_33_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_34_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_35_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_36_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_37_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_38_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_39_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_40_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_206 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_41_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_208 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_42_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_216 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_43_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_218 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_44_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_45_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_226 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_46_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_47_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_234 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_48_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_49_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_238 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_50_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_246 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_51_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_248 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_52_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_53_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_254 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_54_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_256 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_55_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_266 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_56_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_57_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_270 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_58_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_272 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_59_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_274 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_60_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_286 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_61_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_290 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_62_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_63_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_310 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_64_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_322 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_65_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_342 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_66_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_344 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_67_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_348 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size4_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_68_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_360 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_69_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_362 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_70_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_364 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_71_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_366 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_72_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_368 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_73_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_378 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_74_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_380 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_75_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_382 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_76_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_386 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_77_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_388 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_78_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_396 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_79_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_398 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_80_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_400 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_81_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_406 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_82_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_408 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_83_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_414 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_84_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_416 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_85_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_418 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_86_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_426 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_87_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_428 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_88_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__4_ -----

//----- Default net type -----
`default_nettype wire



