//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[2][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Oct 17 11:38:19 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_2__4_ -----
module sb_2__4_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:159] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:159] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:159] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_;
//----- INPUT PORTS -----
input [0:159] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:159] chany_top_out;
//----- OUTPUT PORTS -----
output [0:159] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:159] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:159] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:7] mux_2level_tapbuf_size10_0_sram;
wire [0:7] mux_2level_tapbuf_size10_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size10_mem_0_ccff_tail;
wire [0:7] mux_2level_tapbuf_size11_0_sram;
wire [0:7] mux_2level_tapbuf_size11_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_10_sram;
wire [0:7] mux_2level_tapbuf_size11_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_11_sram;
wire [0:7] mux_2level_tapbuf_size11_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_12_sram;
wire [0:7] mux_2level_tapbuf_size11_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_13_sram;
wire [0:7] mux_2level_tapbuf_size11_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_14_sram;
wire [0:7] mux_2level_tapbuf_size11_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_15_sram;
wire [0:7] mux_2level_tapbuf_size11_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_16_sram;
wire [0:7] mux_2level_tapbuf_size11_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_17_sram;
wire [0:7] mux_2level_tapbuf_size11_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_18_sram;
wire [0:7] mux_2level_tapbuf_size11_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_19_sram;
wire [0:7] mux_2level_tapbuf_size11_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_1_sram;
wire [0:7] mux_2level_tapbuf_size11_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_20_sram;
wire [0:7] mux_2level_tapbuf_size11_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_21_sram;
wire [0:7] mux_2level_tapbuf_size11_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_22_sram;
wire [0:7] mux_2level_tapbuf_size11_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_23_sram;
wire [0:7] mux_2level_tapbuf_size11_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_24_sram;
wire [0:7] mux_2level_tapbuf_size11_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_25_sram;
wire [0:7] mux_2level_tapbuf_size11_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_26_sram;
wire [0:7] mux_2level_tapbuf_size11_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_27_sram;
wire [0:7] mux_2level_tapbuf_size11_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_28_sram;
wire [0:7] mux_2level_tapbuf_size11_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_29_sram;
wire [0:7] mux_2level_tapbuf_size11_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_2_sram;
wire [0:7] mux_2level_tapbuf_size11_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_30_sram;
wire [0:7] mux_2level_tapbuf_size11_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_31_sram;
wire [0:7] mux_2level_tapbuf_size11_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_32_sram;
wire [0:7] mux_2level_tapbuf_size11_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_33_sram;
wire [0:7] mux_2level_tapbuf_size11_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_34_sram;
wire [0:7] mux_2level_tapbuf_size11_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_35_sram;
wire [0:7] mux_2level_tapbuf_size11_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_36_sram;
wire [0:7] mux_2level_tapbuf_size11_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_37_sram;
wire [0:7] mux_2level_tapbuf_size11_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_38_sram;
wire [0:7] mux_2level_tapbuf_size11_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_3_sram;
wire [0:7] mux_2level_tapbuf_size11_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_4_sram;
wire [0:7] mux_2level_tapbuf_size11_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_5_sram;
wire [0:7] mux_2level_tapbuf_size11_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_6_sram;
wire [0:7] mux_2level_tapbuf_size11_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_7_sram;
wire [0:7] mux_2level_tapbuf_size11_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_8_sram;
wire [0:7] mux_2level_tapbuf_size11_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size11_9_sram;
wire [0:7] mux_2level_tapbuf_size11_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size11_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size12_0_sram;
wire [0:7] mux_2level_tapbuf_size12_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_10_sram;
wire [0:7] mux_2level_tapbuf_size12_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_11_sram;
wire [0:7] mux_2level_tapbuf_size12_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_12_sram;
wire [0:7] mux_2level_tapbuf_size12_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_13_sram;
wire [0:7] mux_2level_tapbuf_size12_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_14_sram;
wire [0:7] mux_2level_tapbuf_size12_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_15_sram;
wire [0:7] mux_2level_tapbuf_size12_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_16_sram;
wire [0:7] mux_2level_tapbuf_size12_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_17_sram;
wire [0:7] mux_2level_tapbuf_size12_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_18_sram;
wire [0:7] mux_2level_tapbuf_size12_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_19_sram;
wire [0:7] mux_2level_tapbuf_size12_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_1_sram;
wire [0:7] mux_2level_tapbuf_size12_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_20_sram;
wire [0:7] mux_2level_tapbuf_size12_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_21_sram;
wire [0:7] mux_2level_tapbuf_size12_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_22_sram;
wire [0:7] mux_2level_tapbuf_size12_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_23_sram;
wire [0:7] mux_2level_tapbuf_size12_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_24_sram;
wire [0:7] mux_2level_tapbuf_size12_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_25_sram;
wire [0:7] mux_2level_tapbuf_size12_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_26_sram;
wire [0:7] mux_2level_tapbuf_size12_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_27_sram;
wire [0:7] mux_2level_tapbuf_size12_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_28_sram;
wire [0:7] mux_2level_tapbuf_size12_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_29_sram;
wire [0:7] mux_2level_tapbuf_size12_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_2_sram;
wire [0:7] mux_2level_tapbuf_size12_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_30_sram;
wire [0:7] mux_2level_tapbuf_size12_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_3_sram;
wire [0:7] mux_2level_tapbuf_size12_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_4_sram;
wire [0:7] mux_2level_tapbuf_size12_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_5_sram;
wire [0:7] mux_2level_tapbuf_size12_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_6_sram;
wire [0:7] mux_2level_tapbuf_size12_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_7_sram;
wire [0:7] mux_2level_tapbuf_size12_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_8_sram;
wire [0:7] mux_2level_tapbuf_size12_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size12_9_sram;
wire [0:7] mux_2level_tapbuf_size12_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size12_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size13_0_sram;
wire [0:7] mux_2level_tapbuf_size13_0_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_10_sram;
wire [0:7] mux_2level_tapbuf_size13_10_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_11_sram;
wire [0:7] mux_2level_tapbuf_size13_11_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_12_sram;
wire [0:7] mux_2level_tapbuf_size13_12_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_13_sram;
wire [0:7] mux_2level_tapbuf_size13_13_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_14_sram;
wire [0:7] mux_2level_tapbuf_size13_14_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_15_sram;
wire [0:7] mux_2level_tapbuf_size13_15_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_16_sram;
wire [0:7] mux_2level_tapbuf_size13_16_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_17_sram;
wire [0:7] mux_2level_tapbuf_size13_17_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_18_sram;
wire [0:7] mux_2level_tapbuf_size13_18_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_19_sram;
wire [0:7] mux_2level_tapbuf_size13_19_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_1_sram;
wire [0:7] mux_2level_tapbuf_size13_1_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_20_sram;
wire [0:7] mux_2level_tapbuf_size13_20_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_21_sram;
wire [0:7] mux_2level_tapbuf_size13_21_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_22_sram;
wire [0:7] mux_2level_tapbuf_size13_22_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_23_sram;
wire [0:7] mux_2level_tapbuf_size13_23_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_24_sram;
wire [0:7] mux_2level_tapbuf_size13_24_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_25_sram;
wire [0:7] mux_2level_tapbuf_size13_25_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_26_sram;
wire [0:7] mux_2level_tapbuf_size13_26_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_27_sram;
wire [0:7] mux_2level_tapbuf_size13_27_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_28_sram;
wire [0:7] mux_2level_tapbuf_size13_28_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_29_sram;
wire [0:7] mux_2level_tapbuf_size13_29_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_2_sram;
wire [0:7] mux_2level_tapbuf_size13_2_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_30_sram;
wire [0:7] mux_2level_tapbuf_size13_30_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_31_sram;
wire [0:7] mux_2level_tapbuf_size13_31_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_32_sram;
wire [0:7] mux_2level_tapbuf_size13_32_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_33_sram;
wire [0:7] mux_2level_tapbuf_size13_33_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_34_sram;
wire [0:7] mux_2level_tapbuf_size13_34_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_35_sram;
wire [0:7] mux_2level_tapbuf_size13_35_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_36_sram;
wire [0:7] mux_2level_tapbuf_size13_36_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_37_sram;
wire [0:7] mux_2level_tapbuf_size13_37_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_38_sram;
wire [0:7] mux_2level_tapbuf_size13_38_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_39_sram;
wire [0:7] mux_2level_tapbuf_size13_39_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_3_sram;
wire [0:7] mux_2level_tapbuf_size13_3_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_40_sram;
wire [0:7] mux_2level_tapbuf_size13_40_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_41_sram;
wire [0:7] mux_2level_tapbuf_size13_41_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_42_sram;
wire [0:7] mux_2level_tapbuf_size13_42_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_43_sram;
wire [0:7] mux_2level_tapbuf_size13_43_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_44_sram;
wire [0:7] mux_2level_tapbuf_size13_44_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_45_sram;
wire [0:7] mux_2level_tapbuf_size13_45_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_46_sram;
wire [0:7] mux_2level_tapbuf_size13_46_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_47_sram;
wire [0:7] mux_2level_tapbuf_size13_47_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_4_sram;
wire [0:7] mux_2level_tapbuf_size13_4_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_5_sram;
wire [0:7] mux_2level_tapbuf_size13_5_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_6_sram;
wire [0:7] mux_2level_tapbuf_size13_6_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_7_sram;
wire [0:7] mux_2level_tapbuf_size13_7_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_8_sram;
wire [0:7] mux_2level_tapbuf_size13_8_sram_inv;
wire [0:7] mux_2level_tapbuf_size13_9_sram;
wire [0:7] mux_2level_tapbuf_size13_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size13_mem_9_ccff_tail;
wire [0:7] mux_2level_tapbuf_size15_0_sram;
wire [0:7] mux_2level_tapbuf_size15_0_sram_inv;
wire [0:0] mux_2level_tapbuf_size15_mem_0_ccff_tail;
wire [0:11] mux_2level_tapbuf_size28_0_sram;
wire [0:11] mux_2level_tapbuf_size28_0_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_10_sram;
wire [0:11] mux_2level_tapbuf_size28_10_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_11_sram;
wire [0:11] mux_2level_tapbuf_size28_11_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_12_sram;
wire [0:11] mux_2level_tapbuf_size28_12_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_13_sram;
wire [0:11] mux_2level_tapbuf_size28_13_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_14_sram;
wire [0:11] mux_2level_tapbuf_size28_14_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_15_sram;
wire [0:11] mux_2level_tapbuf_size28_15_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_16_sram;
wire [0:11] mux_2level_tapbuf_size28_16_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_17_sram;
wire [0:11] mux_2level_tapbuf_size28_17_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_18_sram;
wire [0:11] mux_2level_tapbuf_size28_18_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_19_sram;
wire [0:11] mux_2level_tapbuf_size28_19_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_1_sram;
wire [0:11] mux_2level_tapbuf_size28_1_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_20_sram;
wire [0:11] mux_2level_tapbuf_size28_20_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_21_sram;
wire [0:11] mux_2level_tapbuf_size28_21_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_22_sram;
wire [0:11] mux_2level_tapbuf_size28_22_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_23_sram;
wire [0:11] mux_2level_tapbuf_size28_23_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_24_sram;
wire [0:11] mux_2level_tapbuf_size28_24_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_25_sram;
wire [0:11] mux_2level_tapbuf_size28_25_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_26_sram;
wire [0:11] mux_2level_tapbuf_size28_26_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_27_sram;
wire [0:11] mux_2level_tapbuf_size28_27_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_28_sram;
wire [0:11] mux_2level_tapbuf_size28_28_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_29_sram;
wire [0:11] mux_2level_tapbuf_size28_29_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_2_sram;
wire [0:11] mux_2level_tapbuf_size28_2_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_30_sram;
wire [0:11] mux_2level_tapbuf_size28_30_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_31_sram;
wire [0:11] mux_2level_tapbuf_size28_31_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_3_sram;
wire [0:11] mux_2level_tapbuf_size28_3_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_4_sram;
wire [0:11] mux_2level_tapbuf_size28_4_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_5_sram;
wire [0:11] mux_2level_tapbuf_size28_5_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_6_sram;
wire [0:11] mux_2level_tapbuf_size28_6_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_7_sram;
wire [0:11] mux_2level_tapbuf_size28_7_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_8_sram;
wire [0:11] mux_2level_tapbuf_size28_8_sram_inv;
wire [0:11] mux_2level_tapbuf_size28_9_sram;
wire [0:11] mux_2level_tapbuf_size28_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size28_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size28_mem_9_ccff_tail;
wire [0:11] mux_2level_tapbuf_size29_0_sram;
wire [0:11] mux_2level_tapbuf_size29_0_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_1_sram;
wire [0:11] mux_2level_tapbuf_size29_1_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_2_sram;
wire [0:11] mux_2level_tapbuf_size29_2_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_3_sram;
wire [0:11] mux_2level_tapbuf_size29_3_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_4_sram;
wire [0:11] mux_2level_tapbuf_size29_4_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_5_sram;
wire [0:11] mux_2level_tapbuf_size29_5_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_6_sram;
wire [0:11] mux_2level_tapbuf_size29_6_sram_inv;
wire [0:11] mux_2level_tapbuf_size29_7_sram;
wire [0:11] mux_2level_tapbuf_size29_7_sram_inv;
wire [0:0] mux_2level_tapbuf_size29_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size29_mem_7_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[1];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[5];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[9];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[13];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[17];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[21];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[25];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[29];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[33];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[37];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[41];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[45];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[49];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[53];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[57];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[61];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[64] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[65];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[68] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[69];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[72] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[73];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[76] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[77];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[80] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[81];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[84] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[85];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[88] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[89];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[92] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[93];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[96] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[97];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[100] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[101];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[104] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[105];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[108] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[109];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[112] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[113];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[116] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[117];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[120] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[121];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[124] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[125];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[128] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[129];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[132] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[133];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[136] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[137];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[140] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[141];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[144] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[145];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[148] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[149];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[152] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[153];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[156] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[157];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[159];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[0] = chanx_right_in[0];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[1];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[3];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[4] = chanx_right_in[4];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[5];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[7];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[8] = chanx_right_in[8];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[9];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[11];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[12] = chanx_right_in[12];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[13];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[15];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[16] = chanx_right_in[16];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[17];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[19];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[20] = chanx_right_in[20];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[21];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[23];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[24] = chanx_right_in[24];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[25];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[27];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[28] = chanx_right_in[28];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[29];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[31];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[64] = chanx_right_in[64];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[65] = chanx_right_in[65];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[67] = chanx_right_in[67];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[68] = chanx_right_in[68];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[69] = chanx_right_in[69];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[71] = chanx_right_in[71];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[72] = chanx_right_in[72];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[73] = chanx_right_in[73];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[75] = chanx_right_in[75];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[76] = chanx_right_in[76];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[77] = chanx_right_in[77];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[79];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[80] = chanx_right_in[80];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[81] = chanx_right_in[81];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[83];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[84] = chanx_right_in[84];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[85];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[87];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[88] = chanx_right_in[88];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[89] = chanx_right_in[89];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[91];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[92] = chanx_right_in[92];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[93] = chanx_right_in[93];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[95];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[96] = chanx_right_in[96];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[97] = chanx_right_in[97];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[99];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[100] = chanx_right_in[100];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[101] = chanx_right_in[101];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[103] = chanx_right_in[103];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[104] = chanx_right_in[104];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[105] = chanx_right_in[105];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[107] = chanx_right_in[107];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[108] = chanx_right_in[108];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[109] = chanx_right_in[109];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[111] = chanx_right_in[111];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[112] = chanx_right_in[112];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[113] = chanx_right_in[113];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[115] = chanx_right_in[115];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[116] = chanx_right_in[116];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[117] = chanx_right_in[117];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[119] = chanx_right_in[119];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[120] = chanx_right_in[120];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[121] = chanx_right_in[121];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[123] = chanx_right_in[123];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[124] = chanx_right_in[124];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[125] = chanx_right_in[125];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[127] = chanx_right_in[127];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[128] = chanx_right_in[128];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[129] = chanx_right_in[129];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[131] = chanx_right_in[131];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[132] = chanx_right_in[132];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[133] = chanx_right_in[133];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[135] = chanx_right_in[135];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[136] = chanx_right_in[136];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[137] = chanx_right_in[137];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[139] = chanx_right_in[139];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[140] = chanx_right_in[140];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[141] = chanx_right_in[141];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[143] = chanx_right_in[143];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[144] = chanx_right_in[144];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[145] = chanx_right_in[145];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[147] = chanx_right_in[147];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[148] = chanx_right_in[148];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[149] = chanx_right_in[149];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[151] = chanx_right_in[151];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[152] = chanx_right_in[152];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[153] = chanx_right_in[153];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[155] = chanx_right_in[155];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[156] = chanx_right_in[156];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[157] = chanx_right_in[157];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[159] = chanx_right_in[159];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[1];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[5];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[9];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[13];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[17];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[21];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[25];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[29];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[33];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[37];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[41];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[45];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[49];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[53];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[57];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[61];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[64];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[65];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[67];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[68];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[69];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[71];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chany_bottom_in[72];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[73];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[75];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chany_bottom_in[76];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[77];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[79];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chany_bottom_in[80];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[81];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[83];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chany_bottom_in[84];
// ----- Local connection due to Wire 425 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[85];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[87];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chany_bottom_in[88];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[89];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[91];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chany_bottom_in[92];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[93];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[95];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[96] = chany_bottom_in[96];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[97];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[99];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[100] = chany_bottom_in[100];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[101];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[103];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[104] = chany_bottom_in[104];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[105];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[107];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[108] = chany_bottom_in[108];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[109];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[111];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[112] = chany_bottom_in[112];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[113];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[115];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chany_bottom_in[116];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[117];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[119];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[120] = chany_bottom_in[120];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[121];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[123];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[124] = chany_bottom_in[124];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[125];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[127];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[128] = chany_bottom_in[128];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[129];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[131];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chany_bottom_in[132];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[133];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[135];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[136] = chany_bottom_in[136];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[137];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[139];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[140] = chany_bottom_in[140];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[141];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[143];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[144] = chany_bottom_in[144];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[145];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[147];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[148] = chany_bottom_in[148];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[149];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[151];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chany_bottom_in[152];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[153];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[155];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[156] = chany_bottom_in[156];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[157];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[159];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[0] = chanx_left_in[0];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[1];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[3];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[4] = chanx_left_in[4];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[5];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[7];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[8] = chanx_left_in[8];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[9];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[11];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[12] = chanx_left_in[12];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[13];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[15];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[16] = chanx_left_in[16];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[17];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[19];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[20] = chanx_left_in[20];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[21];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[23];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[24] = chanx_left_in[24];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[25];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[27];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[28] = chanx_left_in[28];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[29];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[31];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[33];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[37];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[41];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[45];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[49];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[53];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[57];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[61];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[64] = chanx_left_in[64];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[65];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[67];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[68] = chanx_left_in[68];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[69];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[71];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[72] = chanx_left_in[72];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[73];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[75];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[76] = chanx_left_in[76];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[77];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[79];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[80] = chanx_left_in[80];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[81];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[83];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[84] = chanx_left_in[84];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[85];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[87];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[88] = chanx_left_in[88];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[89];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[91];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[92] = chanx_left_in[92];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[93];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[95];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[96] = chanx_left_in[96];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[97];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[99];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[100] = chanx_left_in[100];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[101];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[103];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[104] = chanx_left_in[104];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[105];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[107];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[108] = chanx_left_in[108];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[109];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[111];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[112] = chanx_left_in[112];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[113];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[115];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[116] = chanx_left_in[116];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[117];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[119];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[120] = chanx_left_in[120];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[121];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[123];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[124] = chanx_left_in[124];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[125];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[127];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[128] = chanx_left_in[128];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[129];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[131];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[132] = chanx_left_in[132];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[133];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[135];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[136] = chanx_left_in[136];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[137];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[139];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[140] = chanx_left_in[140];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[141];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[143];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[144] = chanx_left_in[144];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[145];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[147];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[148] = chanx_left_in[148];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[149];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[151];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[152] = chanx_left_in[152];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[153];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[155];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[156] = chanx_left_in[156];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[157];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[159];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size13 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[1], chanx_right_in[6], chanx_right_in[55], chanx_right_in[108], chany_bottom_in[2], chanx_left_in[0], chanx_left_in[2], chanx_left_in[53], chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size13_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_0_sram_inv[0:7]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size13 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[3], chanx_right_in[10], chanx_right_in[56], chanx_right_in[109], chany_bottom_in[6], chanx_left_in[52], chanx_left_in[105], chanx_left_in[158:159]}),
		.sram(mux_2level_tapbuf_size13_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_1_sram_inv[0:7]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size13 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[4], chanx_right_in[14], chanx_right_in[57], chanx_right_in[111], chany_bottom_in[10], chanx_left_in[51], chanx_left_in[104], chanx_left_in[154], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size13_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_2_sram_inv[0:7]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size13 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[5], chanx_right_in[18], chanx_right_in[59], chanx_right_in[112], chany_bottom_in[14], chanx_left_in[49], chanx_left_in[103], chanx_left_in[150], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size13_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_3_sram_inv[0:7]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size13 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[7], chanx_right_in[22], chanx_right_in[60], chanx_right_in[113], chany_bottom_in[18], chanx_left_in[48], chanx_left_in[101], chanx_left_in[146], chanx_left_in[155]}),
		.sram(mux_2level_tapbuf_size13_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_4_sram_inv[0:7]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size13 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[8], chanx_right_in[26], chanx_right_in[61], chanx_right_in[115], chany_bottom_in[22], chanx_left_in[47], chanx_left_in[100], chanx_left_in[142], chanx_left_in[153]}),
		.sram(mux_2level_tapbuf_size13_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_5_sram_inv[0:7]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size13 mux_top_track_52 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[9], chanx_right_in[30], chanx_right_in[63], chanx_right_in[116], chany_bottom_in[26], chanx_left_in[45], chanx_left_in[99], chanx_left_in[138], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size13_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_6_sram_inv[0:7]),
		.out(chany_top_out[26]));

	mux_2level_tapbuf_size13 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[11], chanx_right_in[34], chanx_right_in[64], chanx_right_in[117], chany_bottom_in[30], chanx_left_in[44], chanx_left_in[97], chanx_left_in[134], chanx_left_in[151]}),
		.sram(mux_2level_tapbuf_size13_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_7_sram_inv[0:7]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size13 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[12], chanx_right_in[38], chanx_right_in[65], chanx_right_in[119], chany_bottom_in[34], chanx_left_in[43], chanx_left_in[96], chanx_left_in[130], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size13_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_8_sram_inv[0:7]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size13 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[13], chanx_right_in[42], chanx_right_in[67], chanx_right_in[120], chany_bottom_in[38], chanx_left_in[41], chanx_left_in[95], chanx_left_in[126], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size13_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_9_sram_inv[0:7]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size13 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[15], chanx_right_in[46], chanx_right_in[68], chanx_right_in[121], chany_bottom_in[42], chanx_left_in[40], chanx_left_in[93], chanx_left_in[122], chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size13_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_10_sram_inv[0:7]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size13 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[16], chanx_right_in[50], chanx_right_in[69], chanx_right_in[123], chany_bottom_in[46], chanx_left_in[39], chanx_left_in[92], chanx_left_in[118], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size13_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_11_sram_inv[0:7]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size13 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[17], chanx_right_in[54], chanx_right_in[71], chanx_right_in[124], chany_bottom_in[50], chanx_left_in[37], chanx_left_in[91], chanx_left_in[114], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size13_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_12_sram_inv[0:7]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size13 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[19], chanx_right_in[58], chanx_right_in[72], chanx_right_in[125], chany_bottom_in[54], chanx_left_in[36], chanx_left_in[89], chanx_left_in[110], chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size13_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_13_sram_inv[0:7]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size13 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[20], chanx_right_in[62], chanx_right_in[73], chanx_right_in[127], chany_bottom_in[58], chanx_left_in[35], chanx_left_in[88], chanx_left_in[106], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size13_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_14_sram_inv[0:7]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size13 mux_top_track_124 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[21], chanx_right_in[66], chanx_right_in[75], chanx_right_in[128], chany_bottom_in[62], chanx_left_in[33], chanx_left_in[87], chanx_left_in[102], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size13_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_15_sram_inv[0:7]),
		.out(chany_top_out[62]));

	mux_2level_tapbuf_size13 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[23], chanx_right_in[70], chanx_right_in[76], chanx_right_in[129], chany_bottom_in[66], chanx_left_in[32], chanx_left_in[85], chanx_left_in[98], chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size13_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_16_sram_inv[0:7]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size13 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[24], chanx_right_in[74], chanx_right_in[77], chanx_right_in[131], chany_bottom_in[70], chanx_left_in[31], chanx_left_in[84], chanx_left_in[94], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size13_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_17_sram_inv[0:7]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size13 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[25], chanx_right_in[78:79], chanx_right_in[132], chany_bottom_in[74], chanx_left_in[29], chanx_left_in[83], chanx_left_in[90], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size13_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_18_sram_inv[0:7]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size13 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[27], chanx_right_in[80], chanx_right_in[82], chanx_right_in[133], chany_bottom_in[78], chanx_left_in[28], chanx_left_in[81], chanx_left_in[86], chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size13_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_19_sram_inv[0:7]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size13 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[28], chanx_right_in[81], chanx_right_in[86], chanx_right_in[135], chany_bottom_in[82], chanx_left_in[27], chanx_left_in[80], chanx_left_in[82], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size13_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_20_sram_inv[0:7]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size13 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[29], chanx_right_in[83], chanx_right_in[90], chanx_right_in[136], chany_bottom_in[86], chanx_left_in[25], chanx_left_in[78:79], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size13_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_21_sram_inv[0:7]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size13 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[31], chanx_right_in[84], chanx_right_in[94], chanx_right_in[137], chany_bottom_in[90], chanx_left_in[24], chanx_left_in[74], chanx_left_in[77], chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size13_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_22_sram_inv[0:7]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size13 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, chanx_right_in[32], chanx_right_in[85], chanx_right_in[98], chanx_right_in[139], chany_bottom_in[94], chanx_left_in[23], chanx_left_in[70], chanx_left_in[76], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size13_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_23_sram_inv[0:7]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size13 mux_top_track_196 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[33], chanx_right_in[87], chanx_right_in[102], chanx_right_in[140], chany_bottom_in[98], chanx_left_in[21], chanx_left_in[66], chanx_left_in[75], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size13_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_24_sram_inv[0:7]),
		.out(chany_top_out[98]));

	mux_2level_tapbuf_size13 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[35], chanx_right_in[88], chanx_right_in[106], chanx_right_in[141], chany_bottom_in[102], chanx_left_in[20], chanx_left_in[62], chanx_left_in[73], chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size13_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_25_sram_inv[0:7]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size13 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[36], chanx_right_in[89], chanx_right_in[110], chanx_right_in[143], chany_bottom_in[106], chanx_left_in[19], chanx_left_in[58], chanx_left_in[72], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size13_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_26_sram_inv[0:7]),
		.out(chany_top_out[106]));

	mux_2level_tapbuf_size13 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[37], chanx_right_in[91], chanx_right_in[114], chanx_right_in[144], chany_bottom_in[110], chanx_left_in[17], chanx_left_in[54], chanx_left_in[71], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size13_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_27_sram_inv[0:7]),
		.out(chany_top_out[110]));

	mux_2level_tapbuf_size13 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[39], chanx_right_in[92], chanx_right_in[118], chanx_right_in[145], chany_bottom_in[114], chanx_left_in[16], chanx_left_in[50], chanx_left_in[69], chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size13_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_28_sram_inv[0:7]),
		.out(chany_top_out[114]));

	mux_2level_tapbuf_size13 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[40], chanx_right_in[93], chanx_right_in[122], chanx_right_in[147], chany_bottom_in[118], chanx_left_in[15], chanx_left_in[46], chanx_left_in[68], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size13_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_29_sram_inv[0:7]),
		.out(chany_top_out[118]));

	mux_2level_tapbuf_size13 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[41], chanx_right_in[95], chanx_right_in[126], chanx_right_in[148], chany_bottom_in[122], chanx_left_in[13], chanx_left_in[42], chanx_left_in[67], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size13_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_30_sram_inv[0:7]),
		.out(chany_top_out[122]));

	mux_2level_tapbuf_size13 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[43], chanx_right_in[96], chanx_right_in[130], chanx_right_in[149], chany_bottom_in[126], chanx_left_in[12], chanx_left_in[38], chanx_left_in[65], chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size13_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_31_sram_inv[0:7]),
		.out(chany_top_out[126]));

	mux_2level_tapbuf_size13 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[44], chanx_right_in[97], chanx_right_in[134], chanx_right_in[151], chany_bottom_in[130], chanx_left_in[11], chanx_left_in[34], chanx_left_in[64], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size13_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_32_sram_inv[0:7]),
		.out(chany_top_out[130]));

	mux_2level_tapbuf_size13 mux_top_track_268 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[45], chanx_right_in[99], chanx_right_in[138], chanx_right_in[152], chany_bottom_in[134], chanx_left_in[9], chanx_left_in[30], chanx_left_in[63], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size13_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_33_sram_inv[0:7]),
		.out(chany_top_out[134]));

	mux_2level_tapbuf_size13 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[47], chanx_right_in[100], chanx_right_in[142], chanx_right_in[153], chany_bottom_in[138], chanx_left_in[8], chanx_left_in[26], chanx_left_in[61], chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size13_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_34_sram_inv[0:7]),
		.out(chany_top_out[138]));

	mux_2level_tapbuf_size13 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[48], chanx_right_in[101], chanx_right_in[146], chanx_right_in[155], chany_bottom_in[142], chanx_left_in[7], chanx_left_in[22], chanx_left_in[60], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size13_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_35_sram_inv[0:7]),
		.out(chany_top_out[142]));

	mux_2level_tapbuf_size13 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[49], chanx_right_in[103], chanx_right_in[150], chanx_right_in[156], chany_bottom_in[146], chanx_left_in[5], chanx_left_in[18], chanx_left_in[59], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size13_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_36_sram_inv[0:7]),
		.out(chany_top_out[146]));

	mux_2level_tapbuf_size13 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[51], chanx_right_in[104], chanx_right_in[154], chanx_right_in[157], chany_bottom_in[150], chanx_left_in[4], chanx_left_in[14], chanx_left_in[57], chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size13_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_37_sram_inv[0:7]),
		.out(chany_top_out[150]));

	mux_2level_tapbuf_size13 mux_top_track_308 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[52], chanx_right_in[105], chanx_right_in[158:159], chany_bottom_in[154], chanx_left_in[3], chanx_left_in[10], chanx_left_in[56], chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size13_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_38_sram_inv[0:7]),
		.out(chany_top_out[154]));

	mux_2level_tapbuf_size13 mux_top_track_316 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, chanx_right_in[0], chanx_right_in[2], chanx_right_in[53], chanx_right_in[107], chany_bottom_in[158], chanx_left_in[1], chanx_left_in[6], chanx_left_in[55], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size13_39_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_39_sram_inv[0:7]),
		.out(chany_top_out[158]));

	mux_2level_tapbuf_size13 mux_right_track_4 (
		.in({chany_top_in[52], chany_top_in[105], chany_top_in[158:159], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[51], chany_bottom_in[104], chany_bottom_in[154], chany_bottom_in[157], chanx_left_in[2]}),
		.sram(mux_2level_tapbuf_size13_40_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_40_sram_inv[0:7]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size13 mux_bottom_track_13 (
		.in({chany_top_in[6], chanx_right_in[49], chanx_right_in[150], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[3], chanx_left_in[10], chanx_left_in[56], chanx_left_in[109]}),
		.sram(mux_2level_tapbuf_size13_41_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_41_sram_inv[0:7]),
		.out(chany_bottom_out[6]));

	mux_2level_tapbuf_size13 mux_bottom_track_21 (
		.in({chany_top_in[10], chanx_right_in[48], chanx_right_in[146], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[4], chanx_left_in[14], chanx_left_in[57], chanx_left_in[111]}),
		.sram(mux_2level_tapbuf_size13_42_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_42_sram_inv[0:7]),
		.out(chany_bottom_out[10]));

	mux_2level_tapbuf_size13 mux_bottom_track_29 (
		.in({chany_top_in[14], chanx_right_in[47], chanx_right_in[142], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[5], chanx_left_in[18], chanx_left_in[59], chanx_left_in[112]}),
		.sram(mux_2level_tapbuf_size13_43_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_43_sram_inv[0:7]),
		.out(chany_bottom_out[14]));

	mux_2level_tapbuf_size13 mux_bottom_track_37 (
		.in({chany_top_in[18], chanx_right_in[45], chanx_right_in[138], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[7], chanx_left_in[22], chanx_left_in[60], chanx_left_in[113]}),
		.sram(mux_2level_tapbuf_size13_44_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_44_sram_inv[0:7]),
		.out(chany_bottom_out[18]));

	mux_2level_tapbuf_size13 mux_bottom_track_45 (
		.in({chany_top_in[22], chanx_right_in[44], chanx_right_in[134], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[8], chanx_left_in[26], chanx_left_in[61], chanx_left_in[115]}),
		.sram(mux_2level_tapbuf_size13_45_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_45_sram_inv[0:7]),
		.out(chany_bottom_out[22]));

	mux_2level_tapbuf_size13 mux_bottom_track_53 (
		.in({chany_top_in[26], chanx_right_in[43], chanx_right_in[130], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[9], chanx_left_in[30], chanx_left_in[63], chanx_left_in[116]}),
		.sram(mux_2level_tapbuf_size13_46_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_46_sram_inv[0:7]),
		.out(chany_bottom_out[26]));

	mux_2level_tapbuf_size13 mux_bottom_track_61 (
		.in({chany_top_in[30], chanx_right_in[41], chanx_right_in[126], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[11], chanx_left_in[34], chanx_left_in[64], chanx_left_in[117]}),
		.sram(mux_2level_tapbuf_size13_47_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size13_47_sram_inv[0:7]),
		.out(chany_bottom_out[30]));

	mux_2level_tapbuf_size13_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_0_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_1_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_2_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_3_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_4_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_5_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_6_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_7_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_8_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_9_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_10_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_11_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_12_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_13_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_14_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_15_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_16_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_17_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_18_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_19_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_20_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_21_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_22_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_23_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_24_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_25_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_26_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_27_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_28_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_29_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_30_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_31_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_32_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_33_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_34_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_35_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_36_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_37_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_38_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_top_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_39_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_39_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_40_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_40_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_41_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_41_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_42_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_42_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_43_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_43_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_37 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_44_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_44_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_45_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_45_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_46_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_46_sram_inv[0:7]));

	mux_2level_tapbuf_size13_mem mem_bottom_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size13_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size13_47_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size13_47_sram_inv[0:7]));

	mux_2level_tapbuf_size11 mux_right_track_12 (
		.in({chany_top_in[0], chany_top_in[2], chany_top_in[53], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[49], chany_bottom_in[150], chanx_left_in[6]}),
		.sram(mux_2level_tapbuf_size11_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_0_sram_inv[0:7]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size11 mux_right_track_20 (
		.in({chany_top_in[1], chany_top_in[6], chany_top_in[55], chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[48], chany_bottom_in[146], chanx_left_in[10]}),
		.sram(mux_2level_tapbuf_size11_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_1_sram_inv[0:7]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size11 mux_right_track_28 (
		.in({chany_top_in[3], chany_top_in[10], chany_top_in[56], chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[47], chany_bottom_in[142], chanx_left_in[14]}),
		.sram(mux_2level_tapbuf_size11_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_2_sram_inv[0:7]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size11 mux_right_track_36 (
		.in({chany_top_in[4], chany_top_in[14], chany_top_in[57], chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[45], chany_bottom_in[138], chanx_left_in[18]}),
		.sram(mux_2level_tapbuf_size11_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_3_sram_inv[0:7]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size11 mux_right_track_44 (
		.in({chany_top_in[5], chany_top_in[18], chany_top_in[59], chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[44], chany_bottom_in[134], chanx_left_in[22]}),
		.sram(mux_2level_tapbuf_size11_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_4_sram_inv[0:7]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size11 mux_right_track_52 (
		.in({chany_top_in[7], chany_top_in[22], chany_top_in[60], chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[43], chany_bottom_in[130], chanx_left_in[26]}),
		.sram(mux_2level_tapbuf_size11_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_5_sram_inv[0:7]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size11 mux_right_track_60 (
		.in({chany_top_in[8], chany_top_in[26], chany_top_in[61], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[41], chany_bottom_in[126], chanx_left_in[30]}),
		.sram(mux_2level_tapbuf_size11_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_6_sram_inv[0:7]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size11 mux_right_track_68 (
		.in({chany_top_in[9], chany_top_in[30], chany_top_in[63], chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[40], chany_bottom_in[122], chanx_left_in[34]}),
		.sram(mux_2level_tapbuf_size11_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_7_sram_inv[0:7]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size11 mux_right_track_76 (
		.in({chany_top_in[11], chany_top_in[34], chany_top_in[64], chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[39], chany_bottom_in[118], chanx_left_in[38]}),
		.sram(mux_2level_tapbuf_size11_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_8_sram_inv[0:7]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size11 mux_right_track_84 (
		.in({chany_top_in[12], chany_top_in[38], chany_top_in[65], chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[37], chany_bottom_in[114], chanx_left_in[42]}),
		.sram(mux_2level_tapbuf_size11_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_9_sram_inv[0:7]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size11 mux_right_track_92 (
		.in({chany_top_in[13], chany_top_in[42], chany_top_in[67], chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[36], chany_bottom_in[110], chanx_left_in[46]}),
		.sram(mux_2level_tapbuf_size11_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_10_sram_inv[0:7]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size11 mux_right_track_100 (
		.in({chany_top_in[15], chany_top_in[46], chany_top_in[68], chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[35], chany_bottom_in[106], chanx_left_in[50]}),
		.sram(mux_2level_tapbuf_size11_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_11_sram_inv[0:7]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size11 mux_right_track_108 (
		.in({chany_top_in[16], chany_top_in[50], chany_top_in[69], chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[33], chany_bottom_in[102], chanx_left_in[54]}),
		.sram(mux_2level_tapbuf_size11_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_12_sram_inv[0:7]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size11 mux_right_track_116 (
		.in({chany_top_in[17], chany_top_in[54], chany_top_in[71], chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[32], chany_bottom_in[98], chanx_left_in[58]}),
		.sram(mux_2level_tapbuf_size11_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_13_sram_inv[0:7]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size11 mux_right_track_124 (
		.in({chany_top_in[19], chany_top_in[58], chany_top_in[72], chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[31], chany_bottom_in[94], chanx_left_in[62]}),
		.sram(mux_2level_tapbuf_size11_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_14_sram_inv[0:7]),
		.out(chanx_right_out[62]));

	mux_2level_tapbuf_size11 mux_right_track_132 (
		.in({chany_top_in[20], chany_top_in[62], chany_top_in[73], chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[29], chany_bottom_in[90], chanx_left_in[66]}),
		.sram(mux_2level_tapbuf_size11_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_15_sram_inv[0:7]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size11 mux_right_track_140 (
		.in({chany_top_in[21], chany_top_in[66], chany_top_in[75], chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[28], chany_bottom_in[86], chanx_left_in[70]}),
		.sram(mux_2level_tapbuf_size11_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_16_sram_inv[0:7]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size11 mux_right_track_148 (
		.in({chany_top_in[23], chany_top_in[70], chany_top_in[76], chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[27], chany_bottom_in[82], chanx_left_in[74]}),
		.sram(mux_2level_tapbuf_size11_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_17_sram_inv[0:7]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size11 mux_right_track_156 (
		.in({chany_top_in[24], chany_top_in[74], chany_top_in[77], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[25], chany_bottom_in[78], chanx_left_in[78]}),
		.sram(mux_2level_tapbuf_size11_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_18_sram_inv[0:7]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size11 mux_right_track_164 (
		.in({chany_top_in[25], chany_top_in[78:79], chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[24], chany_bottom_in[74], chanx_left_in[82]}),
		.sram(mux_2level_tapbuf_size11_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_19_sram_inv[0:7]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size11 mux_right_track_172 (
		.in({chany_top_in[27], chany_top_in[80], chany_top_in[82], chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[23], chany_bottom_in[70], chanx_left_in[86]}),
		.sram(mux_2level_tapbuf_size11_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_20_sram_inv[0:7]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size11 mux_right_track_180 (
		.in({chany_top_in[28], chany_top_in[81], chany_top_in[86], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[21], chany_bottom_in[66], chanx_left_in[90]}),
		.sram(mux_2level_tapbuf_size11_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_21_sram_inv[0:7]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size11 mux_right_track_188 (
		.in({chany_top_in[29], chany_top_in[83], chany_top_in[90], chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[20], chany_bottom_in[62], chanx_left_in[94]}),
		.sram(mux_2level_tapbuf_size11_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_22_sram_inv[0:7]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size11 mux_right_track_196 (
		.in({chany_top_in[31], chany_top_in[84], chany_top_in[94], chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[19], chany_bottom_in[58], chanx_left_in[98]}),
		.sram(mux_2level_tapbuf_size11_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_23_sram_inv[0:7]),
		.out(chanx_right_out[98]));

	mux_2level_tapbuf_size11 mux_right_track_204 (
		.in({chany_top_in[32], chany_top_in[85], chany_top_in[98], chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[17], chany_bottom_in[54], chanx_left_in[102]}),
		.sram(mux_2level_tapbuf_size11_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_24_sram_inv[0:7]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size11 mux_right_track_212 (
		.in({chany_top_in[33], chany_top_in[87], chany_top_in[102], chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[16], chany_bottom_in[50], chanx_left_in[106]}),
		.sram(mux_2level_tapbuf_size11_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_25_sram_inv[0:7]),
		.out(chanx_right_out[106]));

	mux_2level_tapbuf_size11 mux_right_track_220 (
		.in({chany_top_in[35], chany_top_in[88], chany_top_in[106], chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[15], chany_bottom_in[46], chanx_left_in[110]}),
		.sram(mux_2level_tapbuf_size11_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_26_sram_inv[0:7]),
		.out(chanx_right_out[110]));

	mux_2level_tapbuf_size11 mux_right_track_228 (
		.in({chany_top_in[36], chany_top_in[89], chany_top_in[110], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[13], chany_bottom_in[42], chanx_left_in[114]}),
		.sram(mux_2level_tapbuf_size11_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_27_sram_inv[0:7]),
		.out(chanx_right_out[114]));

	mux_2level_tapbuf_size11 mux_right_track_236 (
		.in({chany_top_in[37], chany_top_in[91], chany_top_in[114], chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[12], chany_bottom_in[38], chanx_left_in[118]}),
		.sram(mux_2level_tapbuf_size11_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_28_sram_inv[0:7]),
		.out(chanx_right_out[118]));

	mux_2level_tapbuf_size11 mux_right_track_244 (
		.in({chany_top_in[39], chany_top_in[92], chany_top_in[118], chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[11], chany_bottom_in[34], chanx_left_in[122]}),
		.sram(mux_2level_tapbuf_size11_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_29_sram_inv[0:7]),
		.out(chanx_right_out[122]));

	mux_2level_tapbuf_size11 mux_right_track_252 (
		.in({chany_top_in[40], chany_top_in[93], chany_top_in[122], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[9], chany_bottom_in[30], chanx_left_in[126]}),
		.sram(mux_2level_tapbuf_size11_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_30_sram_inv[0:7]),
		.out(chanx_right_out[126]));

	mux_2level_tapbuf_size11 mux_right_track_260 (
		.in({chany_top_in[41], chany_top_in[95], chany_top_in[126], chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[8], chany_bottom_in[26], chanx_left_in[130]}),
		.sram(mux_2level_tapbuf_size11_31_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_31_sram_inv[0:7]),
		.out(chanx_right_out[130]));

	mux_2level_tapbuf_size11 mux_right_track_268 (
		.in({chany_top_in[43], chany_top_in[96], chany_top_in[130], chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[7], chany_bottom_in[22], chanx_left_in[134]}),
		.sram(mux_2level_tapbuf_size11_32_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_32_sram_inv[0:7]),
		.out(chanx_right_out[134]));

	mux_2level_tapbuf_size11 mux_right_track_276 (
		.in({chany_top_in[44], chany_top_in[97], chany_top_in[134], chany_top_in[151], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[5], chany_bottom_in[18], chanx_left_in[138]}),
		.sram(mux_2level_tapbuf_size11_33_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_33_sram_inv[0:7]),
		.out(chanx_right_out[138]));

	mux_2level_tapbuf_size11 mux_right_track_284 (
		.in({chany_top_in[45], chany_top_in[99], chany_top_in[138], chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[4], chany_bottom_in[14], chanx_left_in[142]}),
		.sram(mux_2level_tapbuf_size11_34_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_34_sram_inv[0:7]),
		.out(chanx_right_out[142]));

	mux_2level_tapbuf_size11 mux_right_track_292 (
		.in({chany_top_in[47], chany_top_in[100], chany_top_in[142], chany_top_in[153], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[3], chany_bottom_in[10], chanx_left_in[146]}),
		.sram(mux_2level_tapbuf_size11_35_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_35_sram_inv[0:7]),
		.out(chanx_right_out[146]));

	mux_2level_tapbuf_size11 mux_right_track_300 (
		.in({chany_top_in[48], chany_top_in[101], chany_top_in[146], chany_top_in[155], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[1], chany_bottom_in[6], chanx_left_in[150]}),
		.sram(mux_2level_tapbuf_size11_36_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_36_sram_inv[0:7]),
		.out(chanx_right_out[150]));

	mux_2level_tapbuf_size11 mux_right_track_308 (
		.in({chany_top_in[49], chany_top_in[103], chany_top_in[150], chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[0], chany_bottom_in[2], chanx_left_in[154]}),
		.sram(mux_2level_tapbuf_size11_37_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_37_sram_inv[0:7]),
		.out(chanx_right_out[154]));

	mux_2level_tapbuf_size11 mux_bottom_track_317 (
		.in({chany_top_in[158], chanx_right_in[158], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[0], chanx_left_in[2], chanx_left_in[53], chanx_left_in[107]}),
		.sram(mux_2level_tapbuf_size11_38_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size11_38_sram_inv[0:7]),
		.out(chany_bottom_out[158]));

	mux_2level_tapbuf_size11_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_0_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_1_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_2_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_3_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_4_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_5_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_6_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_7_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_8_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_9_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_10_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_11_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_12_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_13_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_124 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_14_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_15_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_16_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_17_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_18_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_19_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_20_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_21_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_22_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_196 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_23_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_24_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_212 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_25_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_220 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_26_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_228 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_27_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_236 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_28_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_244 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_29_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_252 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_30_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_260 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_31_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_31_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_268 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_32_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_32_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_276 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_33_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_33_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_284 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_34_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_34_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_292 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_35_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_35_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_300 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_36_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_36_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_right_track_308 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_37_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_37_sram_inv[0:7]));

	mux_2level_tapbuf_size11_mem mem_bottom_track_317 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size11_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size11_38_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size11_38_sram_inv[0:7]));

	mux_2level_tapbuf_size10 mux_right_track_316 (
		.in({chany_top_in[51], chany_top_in[104], chany_top_in[154], chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[158], chanx_left_in[158]}),
		.sram(mux_2level_tapbuf_size10_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size10_0_sram_inv[0:7]),
		.out(chanx_right_out[158]));

	mux_2level_tapbuf_size10_mem mem_right_track_316 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size10_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size10_0_sram_inv[0:7]));

	mux_2level_tapbuf_size15 mux_bottom_track_5 (
		.in({chany_top_in[2], chanx_right_in[51], chanx_right_in[104], chanx_right_in[154], chanx_right_in[157], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[1], chanx_left_in[6], chanx_left_in[55], chanx_left_in[108]}),
		.sram(mux_2level_tapbuf_size15_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size15_0_sram_inv[0:7]),
		.out(chany_bottom_out[2]));

	mux_2level_tapbuf_size15_mem mem_bottom_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size15_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size15_0_sram_inv[0:7]));

	mux_2level_tapbuf_size12 mux_bottom_track_69 (
		.in({chany_top_in[34], chanx_right_in[40], chanx_right_in[122], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[12], chanx_left_in[38], chanx_left_in[65], chanx_left_in[119]}),
		.sram(mux_2level_tapbuf_size12_0_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_0_sram_inv[0:7]),
		.out(chany_bottom_out[34]));

	mux_2level_tapbuf_size12 mux_bottom_track_77 (
		.in({chany_top_in[38], chanx_right_in[39], chanx_right_in[118], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[13], chanx_left_in[42], chanx_left_in[67], chanx_left_in[120]}),
		.sram(mux_2level_tapbuf_size12_1_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_1_sram_inv[0:7]),
		.out(chany_bottom_out[38]));

	mux_2level_tapbuf_size12 mux_bottom_track_85 (
		.in({chany_top_in[42], chanx_right_in[37], chanx_right_in[114], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[15], chanx_left_in[46], chanx_left_in[68], chanx_left_in[121]}),
		.sram(mux_2level_tapbuf_size12_2_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_2_sram_inv[0:7]),
		.out(chany_bottom_out[42]));

	mux_2level_tapbuf_size12 mux_bottom_track_93 (
		.in({chany_top_in[46], chanx_right_in[36], chanx_right_in[110], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[16], chanx_left_in[50], chanx_left_in[69], chanx_left_in[123]}),
		.sram(mux_2level_tapbuf_size12_3_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_3_sram_inv[0:7]),
		.out(chany_bottom_out[46]));

	mux_2level_tapbuf_size12 mux_bottom_track_101 (
		.in({chany_top_in[50], chanx_right_in[35], chanx_right_in[106], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[17], chanx_left_in[54], chanx_left_in[71], chanx_left_in[124]}),
		.sram(mux_2level_tapbuf_size12_4_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_4_sram_inv[0:7]),
		.out(chany_bottom_out[50]));

	mux_2level_tapbuf_size12 mux_bottom_track_109 (
		.in({chany_top_in[54], chanx_right_in[33], chanx_right_in[102], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[19], chanx_left_in[58], chanx_left_in[72], chanx_left_in[125]}),
		.sram(mux_2level_tapbuf_size12_5_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_5_sram_inv[0:7]),
		.out(chany_bottom_out[54]));

	mux_2level_tapbuf_size12 mux_bottom_track_117 (
		.in({chany_top_in[58], chanx_right_in[32], chanx_right_in[98], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[20], chanx_left_in[62], chanx_left_in[73], chanx_left_in[127]}),
		.sram(mux_2level_tapbuf_size12_6_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_6_sram_inv[0:7]),
		.out(chany_bottom_out[58]));

	mux_2level_tapbuf_size12 mux_bottom_track_125 (
		.in({chany_top_in[62], chanx_right_in[31], chanx_right_in[94], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_1_, chanx_left_in[21], chanx_left_in[66], chanx_left_in[75], chanx_left_in[128]}),
		.sram(mux_2level_tapbuf_size12_7_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_7_sram_inv[0:7]),
		.out(chany_bottom_out[62]));

	mux_2level_tapbuf_size12 mux_bottom_track_133 (
		.in({chany_top_in[66], chanx_right_in[29], chanx_right_in[90], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[23], chanx_left_in[70], chanx_left_in[76], chanx_left_in[129]}),
		.sram(mux_2level_tapbuf_size12_8_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_8_sram_inv[0:7]),
		.out(chany_bottom_out[66]));

	mux_2level_tapbuf_size12 mux_bottom_track_141 (
		.in({chany_top_in[70], chanx_right_in[28], chanx_right_in[86], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[24], chanx_left_in[74], chanx_left_in[77], chanx_left_in[131]}),
		.sram(mux_2level_tapbuf_size12_9_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_9_sram_inv[0:7]),
		.out(chany_bottom_out[70]));

	mux_2level_tapbuf_size12 mux_bottom_track_149 (
		.in({chany_top_in[74], chanx_right_in[27], chanx_right_in[82], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[25], chanx_left_in[78:79], chanx_left_in[132]}),
		.sram(mux_2level_tapbuf_size12_10_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_10_sram_inv[0:7]),
		.out(chany_bottom_out[74]));

	mux_2level_tapbuf_size12 mux_bottom_track_157 (
		.in({chany_top_in[78], chanx_right_in[25], chanx_right_in[78], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[27], chanx_left_in[80], chanx_left_in[82], chanx_left_in[133]}),
		.sram(mux_2level_tapbuf_size12_11_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_11_sram_inv[0:7]),
		.out(chany_bottom_out[78]));

	mux_2level_tapbuf_size12 mux_bottom_track_165 (
		.in({chany_top_in[82], chanx_right_in[24], chanx_right_in[74], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[28], chanx_left_in[81], chanx_left_in[86], chanx_left_in[135]}),
		.sram(mux_2level_tapbuf_size12_12_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_12_sram_inv[0:7]),
		.out(chany_bottom_out[82]));

	mux_2level_tapbuf_size12 mux_bottom_track_173 (
		.in({chany_top_in[86], chanx_right_in[23], chanx_right_in[70], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[29], chanx_left_in[83], chanx_left_in[90], chanx_left_in[136]}),
		.sram(mux_2level_tapbuf_size12_13_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_13_sram_inv[0:7]),
		.out(chany_bottom_out[86]));

	mux_2level_tapbuf_size12 mux_bottom_track_181 (
		.in({chany_top_in[90], chanx_right_in[21], chanx_right_in[66], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[31], chanx_left_in[84], chanx_left_in[94], chanx_left_in[137]}),
		.sram(mux_2level_tapbuf_size12_14_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_14_sram_inv[0:7]),
		.out(chany_bottom_out[90]));

	mux_2level_tapbuf_size12 mux_bottom_track_189 (
		.in({chany_top_in[94], chanx_right_in[20], chanx_right_in[62], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[32], chanx_left_in[85], chanx_left_in[98], chanx_left_in[139]}),
		.sram(mux_2level_tapbuf_size12_15_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_15_sram_inv[0:7]),
		.out(chany_bottom_out[94]));

	mux_2level_tapbuf_size12 mux_bottom_track_197 (
		.in({chany_top_in[98], chanx_right_in[19], chanx_right_in[58], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[33], chanx_left_in[87], chanx_left_in[102], chanx_left_in[140]}),
		.sram(mux_2level_tapbuf_size12_16_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_16_sram_inv[0:7]),
		.out(chany_bottom_out[98]));

	mux_2level_tapbuf_size12 mux_bottom_track_205 (
		.in({chany_top_in[102], chanx_right_in[17], chanx_right_in[54], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[35], chanx_left_in[88], chanx_left_in[106], chanx_left_in[141]}),
		.sram(mux_2level_tapbuf_size12_17_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_17_sram_inv[0:7]),
		.out(chany_bottom_out[102]));

	mux_2level_tapbuf_size12 mux_bottom_track_213 (
		.in({chany_top_in[106], chanx_right_in[16], chanx_right_in[50], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[36], chanx_left_in[89], chanx_left_in[110], chanx_left_in[143]}),
		.sram(mux_2level_tapbuf_size12_18_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_18_sram_inv[0:7]),
		.out(chany_bottom_out[106]));

	mux_2level_tapbuf_size12 mux_bottom_track_221 (
		.in({chany_top_in[110], chanx_right_in[15], chanx_right_in[46], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[37], chanx_left_in[91], chanx_left_in[114], chanx_left_in[144]}),
		.sram(mux_2level_tapbuf_size12_19_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_19_sram_inv[0:7]),
		.out(chany_bottom_out[110]));

	mux_2level_tapbuf_size12 mux_bottom_track_229 (
		.in({chany_top_in[114], chanx_right_in[13], chanx_right_in[42], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[39], chanx_left_in[92], chanx_left_in[118], chanx_left_in[145]}),
		.sram(mux_2level_tapbuf_size12_20_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_20_sram_inv[0:7]),
		.out(chany_bottom_out[114]));

	mux_2level_tapbuf_size12 mux_bottom_track_237 (
		.in({chany_top_in[118], chanx_right_in[12], chanx_right_in[38], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[40], chanx_left_in[93], chanx_left_in[122], chanx_left_in[147]}),
		.sram(mux_2level_tapbuf_size12_21_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_21_sram_inv[0:7]),
		.out(chany_bottom_out[118]));

	mux_2level_tapbuf_size12 mux_bottom_track_245 (
		.in({chany_top_in[122], chanx_right_in[11], chanx_right_in[34], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[41], chanx_left_in[95], chanx_left_in[126], chanx_left_in[148]}),
		.sram(mux_2level_tapbuf_size12_22_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_22_sram_inv[0:7]),
		.out(chany_bottom_out[122]));

	mux_2level_tapbuf_size12 mux_bottom_track_253 (
		.in({chany_top_in[126], chanx_right_in[9], chanx_right_in[30], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_, chanx_left_in[43], chanx_left_in[96], chanx_left_in[130], chanx_left_in[149]}),
		.sram(mux_2level_tapbuf_size12_23_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_23_sram_inv[0:7]),
		.out(chany_bottom_out[126]));

	mux_2level_tapbuf_size12 mux_bottom_track_261 (
		.in({chany_top_in[130], chanx_right_in[8], chanx_right_in[26], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[44], chanx_left_in[97], chanx_left_in[134], chanx_left_in[151]}),
		.sram(mux_2level_tapbuf_size12_24_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_24_sram_inv[0:7]),
		.out(chany_bottom_out[130]));

	mux_2level_tapbuf_size12 mux_bottom_track_269 (
		.in({chany_top_in[134], chanx_right_in[7], chanx_right_in[22], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[45], chanx_left_in[99], chanx_left_in[138], chanx_left_in[152]}),
		.sram(mux_2level_tapbuf_size12_25_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_25_sram_inv[0:7]),
		.out(chany_bottom_out[134]));

	mux_2level_tapbuf_size12 mux_bottom_track_277 (
		.in({chany_top_in[138], chanx_right_in[5], chanx_right_in[18], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[47], chanx_left_in[100], chanx_left_in[142], chanx_left_in[153]}),
		.sram(mux_2level_tapbuf_size12_26_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_26_sram_inv[0:7]),
		.out(chany_bottom_out[138]));

	mux_2level_tapbuf_size12 mux_bottom_track_285 (
		.in({chany_top_in[142], chanx_right_in[4], chanx_right_in[14], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[48], chanx_left_in[101], chanx_left_in[146], chanx_left_in[155]}),
		.sram(mux_2level_tapbuf_size12_27_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_27_sram_inv[0:7]),
		.out(chany_bottom_out[142]));

	mux_2level_tapbuf_size12 mux_bottom_track_293 (
		.in({chany_top_in[146], chanx_right_in[3], chanx_right_in[10], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[49], chanx_left_in[103], chanx_left_in[150], chanx_left_in[156]}),
		.sram(mux_2level_tapbuf_size12_28_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_28_sram_inv[0:7]),
		.out(chany_bottom_out[146]));

	mux_2level_tapbuf_size12 mux_bottom_track_301 (
		.in({chany_top_in[150], chanx_right_in[1], chanx_right_in[6], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[51], chanx_left_in[104], chanx_left_in[154], chanx_left_in[157]}),
		.sram(mux_2level_tapbuf_size12_29_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_29_sram_inv[0:7]),
		.out(chany_bottom_out[150]));

	mux_2level_tapbuf_size12 mux_bottom_track_309 (
		.in({chany_top_in[154], chanx_right_in[0], chanx_right_in[2], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_1_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_1_, chanx_left_in[52], chanx_left_in[105], chanx_left_in[158:159]}),
		.sram(mux_2level_tapbuf_size12_30_sram[0:7]),
		.sram_inv(mux_2level_tapbuf_size12_30_sram_inv[0:7]),
		.out(chany_bottom_out[154]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size13_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_0_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_0_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_77 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_1_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_1_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_2_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_2_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_3_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_3_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_101 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_4_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_4_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_109 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_5_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_5_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_117 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_6_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_6_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_125 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_7_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_7_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_133 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_8_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_8_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_141 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_9_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_9_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_149 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_10_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_10_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_157 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_11_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_11_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_165 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_12_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_12_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_173 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_13_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_13_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_181 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_14_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_14_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_189 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_15_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_15_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_197 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_16_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_16_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_205 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_17_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_17_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_213 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_18_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_18_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_221 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_19_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_19_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_229 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_20_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_20_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_237 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_21_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_21_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_245 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_22_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_22_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_253 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_23_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_23_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_261 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_24_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_24_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_269 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_25_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_25_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_277 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_26_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_26_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_285 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_27_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_27_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_293 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_28_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_28_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_301 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_29_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_29_sram_inv[0:7]));

	mux_2level_tapbuf_size12_mem mem_bottom_track_309 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size12_30_sram[0:7]),
		.mem_outb(mux_2level_tapbuf_size12_30_sram_inv[0:7]));

	mux_2level_tapbuf_size29 mux_left_track_5 (
		.in({chany_top_in[0], chany_top_in[2], chany_top_in[53], chany_top_in[107], chanx_right_in[2], chany_bottom_in[52], chany_bottom_in[105], chany_bottom_in[158:159], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_0_sram_inv[0:11]),
		.out(chanx_left_out[2]));

	mux_2level_tapbuf_size29 mux_left_track_13 (
		.in({chany_top_in[52], chany_top_in[105], chany_top_in[158:159], chanx_right_in[6], chany_bottom_in[0], chany_bottom_in[2], chany_bottom_in[53], chany_bottom_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_1_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_1_sram_inv[0:11]),
		.out(chanx_left_out[6]));

	mux_2level_tapbuf_size29 mux_left_track_21 (
		.in({chany_top_in[51], chany_top_in[104], chany_top_in[154], chany_top_in[157], chanx_right_in[10], chany_bottom_in[1], chany_bottom_in[6], chany_bottom_in[55], chany_bottom_in[108], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_2_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_2_sram_inv[0:11]),
		.out(chanx_left_out[10]));

	mux_2level_tapbuf_size29 mux_left_track_29 (
		.in({chany_top_in[49], chany_top_in[103], chany_top_in[150], chany_top_in[156], chanx_right_in[14], chany_bottom_in[3], chany_bottom_in[10], chany_bottom_in[56], chany_bottom_in[109], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_3_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_3_sram_inv[0:11]),
		.out(chanx_left_out[14]));

	mux_2level_tapbuf_size29 mux_left_track_37 (
		.in({chany_top_in[48], chany_top_in[101], chany_top_in[146], chany_top_in[155], chanx_right_in[18], chany_bottom_in[4], chany_bottom_in[14], chany_bottom_in[57], chany_bottom_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_4_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_4_sram_inv[0:11]),
		.out(chanx_left_out[18]));

	mux_2level_tapbuf_size29 mux_left_track_45 (
		.in({chany_top_in[47], chany_top_in[100], chany_top_in[142], chany_top_in[153], chanx_right_in[22], chany_bottom_in[5], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[112], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_5_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_5_sram_inv[0:11]),
		.out(chanx_left_out[22]));

	mux_2level_tapbuf_size29 mux_left_track_53 (
		.in({chany_top_in[45], chany_top_in[99], chany_top_in[138], chany_top_in[152], chanx_right_in[26], chany_bottom_in[7], chany_bottom_in[22], chany_bottom_in[60], chany_bottom_in[113], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_6_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_6_sram_inv[0:11]),
		.out(chanx_left_out[26]));

	mux_2level_tapbuf_size29 mux_left_track_61 (
		.in({chany_top_in[44], chany_top_in[97], chany_top_in[134], chany_top_in[151], chanx_right_in[30], chany_bottom_in[8], chany_bottom_in[26], chany_bottom_in[61], chany_bottom_in[115], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size29_7_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size29_7_sram_inv[0:11]),
		.out(chanx_left_out[30]));

	mux_2level_tapbuf_size29_mem mem_left_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size11_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_0_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_1_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_1_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_2_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_2_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_3_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_3_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_37 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_4_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_4_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_5_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_5_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_6_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_6_sram_inv[0:11]));

	mux_2level_tapbuf_size29_mem mem_left_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size29_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size29_7_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size29_7_sram_inv[0:11]));

	mux_2level_tapbuf_size28 mux_left_track_69 (
		.in({chany_top_in[43], chany_top_in[96], chany_top_in[130], chany_top_in[149], chanx_right_in[34], chany_bottom_in[9], chany_bottom_in[30], chany_bottom_in[63], chany_bottom_in[116], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_0_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_0_sram_inv[0:11]),
		.out(chanx_left_out[34]));

	mux_2level_tapbuf_size28 mux_left_track_77 (
		.in({chany_top_in[41], chany_top_in[95], chany_top_in[126], chany_top_in[148], chanx_right_in[38], chany_bottom_in[11], chany_bottom_in[34], chany_bottom_in[64], chany_bottom_in[117], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_1_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_1_sram_inv[0:11]),
		.out(chanx_left_out[38]));

	mux_2level_tapbuf_size28 mux_left_track_85 (
		.in({chany_top_in[40], chany_top_in[93], chany_top_in[122], chany_top_in[147], chanx_right_in[42], chany_bottom_in[12], chany_bottom_in[38], chany_bottom_in[65], chany_bottom_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_2_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_2_sram_inv[0:11]),
		.out(chanx_left_out[42]));

	mux_2level_tapbuf_size28 mux_left_track_93 (
		.in({chany_top_in[39], chany_top_in[92], chany_top_in[118], chany_top_in[145], chanx_right_in[46], chany_bottom_in[13], chany_bottom_in[42], chany_bottom_in[67], chany_bottom_in[120], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_3_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_3_sram_inv[0:11]),
		.out(chanx_left_out[46]));

	mux_2level_tapbuf_size28 mux_left_track_101 (
		.in({chany_top_in[37], chany_top_in[91], chany_top_in[114], chany_top_in[144], chanx_right_in[50], chany_bottom_in[15], chany_bottom_in[46], chany_bottom_in[68], chany_bottom_in[121], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_4_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_4_sram_inv[0:11]),
		.out(chanx_left_out[50]));

	mux_2level_tapbuf_size28 mux_left_track_109 (
		.in({chany_top_in[36], chany_top_in[89], chany_top_in[110], chany_top_in[143], chanx_right_in[54], chany_bottom_in[16], chany_bottom_in[50], chany_bottom_in[69], chany_bottom_in[123], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_5_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_5_sram_inv[0:11]),
		.out(chanx_left_out[54]));

	mux_2level_tapbuf_size28 mux_left_track_117 (
		.in({chany_top_in[35], chany_top_in[88], chany_top_in[106], chany_top_in[141], chanx_right_in[58], chany_bottom_in[17], chany_bottom_in[54], chany_bottom_in[71], chany_bottom_in[124], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_6_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_6_sram_inv[0:11]),
		.out(chanx_left_out[58]));

	mux_2level_tapbuf_size28 mux_left_track_125 (
		.in({chany_top_in[33], chany_top_in[87], chany_top_in[102], chany_top_in[140], chanx_right_in[62], chany_bottom_in[19], chany_bottom_in[58], chany_bottom_in[72], chany_bottom_in[125], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_25_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.sram(mux_2level_tapbuf_size28_7_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_7_sram_inv[0:11]),
		.out(chanx_left_out[62]));

	mux_2level_tapbuf_size28 mux_left_track_133 (
		.in({chany_top_in[32], chany_top_in[85], chany_top_in[98], chany_top_in[139], chanx_right_in[66], chany_bottom_in[20], chany_bottom_in[62], chany_bottom_in[73], chany_bottom_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_8_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_8_sram_inv[0:11]),
		.out(chanx_left_out[66]));

	mux_2level_tapbuf_size28 mux_left_track_141 (
		.in({chany_top_in[31], chany_top_in[84], chany_top_in[94], chany_top_in[137], chanx_right_in[70], chany_bottom_in[21], chany_bottom_in[66], chany_bottom_in[75], chany_bottom_in[128], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_9_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_9_sram_inv[0:11]),
		.out(chanx_left_out[70]));

	mux_2level_tapbuf_size28 mux_left_track_149 (
		.in({chany_top_in[29], chany_top_in[83], chany_top_in[90], chany_top_in[136], chanx_right_in[74], chany_bottom_in[23], chany_bottom_in[70], chany_bottom_in[76], chany_bottom_in[129], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_10_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_10_sram_inv[0:11]),
		.out(chanx_left_out[74]));

	mux_2level_tapbuf_size28 mux_left_track_157 (
		.in({chany_top_in[28], chany_top_in[81], chany_top_in[86], chany_top_in[135], chanx_right_in[78], chany_bottom_in[24], chany_bottom_in[74], chany_bottom_in[77], chany_bottom_in[131], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_11_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_11_sram_inv[0:11]),
		.out(chanx_left_out[78]));

	mux_2level_tapbuf_size28 mux_left_track_165 (
		.in({chany_top_in[27], chany_top_in[80], chany_top_in[82], chany_top_in[133], chanx_right_in[82], chany_bottom_in[25], chany_bottom_in[78:79], chany_bottom_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_12_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_12_sram_inv[0:11]),
		.out(chanx_left_out[82]));

	mux_2level_tapbuf_size28 mux_left_track_173 (
		.in({chany_top_in[25], chany_top_in[78:79], chany_top_in[132], chanx_right_in[86], chany_bottom_in[27], chany_bottom_in[80], chany_bottom_in[82], chany_bottom_in[133], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_13_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_13_sram_inv[0:11]),
		.out(chanx_left_out[86]));

	mux_2level_tapbuf_size28 mux_left_track_181 (
		.in({chany_top_in[24], chany_top_in[74], chany_top_in[77], chany_top_in[131], chanx_right_in[90], chany_bottom_in[28], chany_bottom_in[81], chany_bottom_in[86], chany_bottom_in[135], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_14_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_14_sram_inv[0:11]),
		.out(chanx_left_out[90]));

	mux_2level_tapbuf_size28 mux_left_track_189 (
		.in({chany_top_in[23], chany_top_in[70], chany_top_in[76], chany_top_in[129], chanx_right_in[94], chany_bottom_in[29], chany_bottom_in[83], chany_bottom_in[90], chany_bottom_in[136], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_23_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_33_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_15_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_15_sram_inv[0:11]),
		.out(chanx_left_out[94]));

	mux_2level_tapbuf_size28 mux_left_track_197 (
		.in({chany_top_in[21], chany_top_in[66], chany_top_in[75], chany_top_in[128], chanx_right_in[98], chany_bottom_in[31], chany_bottom_in[84], chany_bottom_in[94], chany_bottom_in[137], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_16_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_16_sram_inv[0:11]),
		.out(chanx_left_out[98]));

	mux_2level_tapbuf_size28 mux_left_track_205 (
		.in({chany_top_in[20], chany_top_in[62], chany_top_in[73], chany_top_in[127], chanx_right_in[102], chany_bottom_in[32], chany_bottom_in[85], chany_bottom_in[98], chany_bottom_in[139], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_17_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_17_sram_inv[0:11]),
		.out(chanx_left_out[102]));

	mux_2level_tapbuf_size28 mux_left_track_213 (
		.in({chany_top_in[19], chany_top_in[58], chany_top_in[72], chany_top_in[125], chanx_right_in[106], chany_bottom_in[33], chany_bottom_in[87], chany_bottom_in[102], chany_bottom_in[140], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_18_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_18_sram_inv[0:11]),
		.out(chanx_left_out[106]));

	mux_2level_tapbuf_size28 mux_left_track_221 (
		.in({chany_top_in[17], chany_top_in[54], chany_top_in[71], chany_top_in[124], chanx_right_in[110], chany_bottom_in[35], chany_bottom_in[88], chany_bottom_in[106], chany_bottom_in[141], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_19_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_19_sram_inv[0:11]),
		.out(chanx_left_out[110]));

	mux_2level_tapbuf_size28 mux_left_track_229 (
		.in({chany_top_in[16], chany_top_in[50], chany_top_in[69], chany_top_in[123], chanx_right_in[114], chany_bottom_in[36], chany_bottom_in[89], chany_bottom_in[110], chany_bottom_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_20_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_20_sram_inv[0:11]),
		.out(chanx_left_out[114]));

	mux_2level_tapbuf_size28 mux_left_track_237 (
		.in({chany_top_in[15], chany_top_in[46], chany_top_in[68], chany_top_in[121], chanx_right_in[118], chany_bottom_in[37], chany_bottom_in[91], chany_bottom_in[114], chany_bottom_in[144], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_21_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_21_sram_inv[0:11]),
		.out(chanx_left_out[118]));

	mux_2level_tapbuf_size28 mux_left_track_245 (
		.in({chany_top_in[13], chany_top_in[42], chany_top_in[67], chany_top_in[120], chanx_right_in[122], chany_bottom_in[39], chany_bottom_in[92], chany_bottom_in[118], chany_bottom_in[145], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_22_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_22_sram_inv[0:11]),
		.out(chanx_left_out[122]));

	mux_2level_tapbuf_size28 mux_left_track_253 (
		.in({chany_top_in[12], chany_top_in[38], chany_top_in[65], chany_top_in[119], chanx_right_in[126], chany_bottom_in[40], chany_bottom_in[93], chany_bottom_in[122], chany_bottom_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_11_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_21_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_31_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_0_}),
		.sram(mux_2level_tapbuf_size28_23_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_23_sram_inv[0:11]),
		.out(chanx_left_out[126]));

	mux_2level_tapbuf_size28 mux_left_track_261 (
		.in({chany_top_in[11], chany_top_in[34], chany_top_in[64], chany_top_in[117], chanx_right_in[130], chany_bottom_in[41], chany_bottom_in[95], chany_bottom_in[126], chany_bottom_in[148], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_24_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_24_sram_inv[0:11]),
		.out(chanx_left_out[130]));

	mux_2level_tapbuf_size28 mux_left_track_269 (
		.in({chany_top_in[9], chany_top_in[30], chany_top_in[63], chany_top_in[116], chanx_right_in[134], chany_bottom_in[43], chany_bottom_in[96], chany_bottom_in[130], chany_bottom_in[149], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_25_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_25_sram_inv[0:11]),
		.out(chanx_left_out[134]));

	mux_2level_tapbuf_size28 mux_left_track_277 (
		.in({chany_top_in[8], chany_top_in[26], chany_top_in[61], chany_top_in[115], chanx_right_in[138], chany_bottom_in[44], chany_bottom_in[97], chany_bottom_in[134], chany_bottom_in[151], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_26_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_26_sram_inv[0:11]),
		.out(chanx_left_out[138]));

	mux_2level_tapbuf_size28 mux_left_track_285 (
		.in({chany_top_in[7], chany_top_in[22], chany_top_in[60], chany_top_in[113], chanx_right_in[142], chany_bottom_in[45], chany_bottom_in[99], chany_bottom_in[138], chany_bottom_in[152], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_27_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_27_sram_inv[0:11]),
		.out(chanx_left_out[142]));

	mux_2level_tapbuf_size28 mux_left_track_293 (
		.in({chany_top_in[5], chany_top_in[18], chany_top_in[59], chany_top_in[112], chanx_right_in[146], chany_bottom_in[47], chany_bottom_in[100], chany_bottom_in[142], chany_bottom_in[153], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_28_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_28_sram_inv[0:11]),
		.out(chanx_left_out[146]));

	mux_2level_tapbuf_size28 mux_left_track_301 (
		.in({chany_top_in[4], chany_top_in[14], chany_top_in[57], chany_top_in[111], chanx_right_in[150], chany_bottom_in[48], chany_bottom_in[101], chany_bottom_in[146], chany_bottom_in[155], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_29_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_29_sram_inv[0:11]),
		.out(chanx_left_out[150]));

	mux_2level_tapbuf_size28 mux_left_track_309 (
		.in({chany_top_in[3], chany_top_in[10], chany_top_in[56], chany_top_in[109], chanx_right_in[154], chany_bottom_in[49], chany_bottom_in[103], chany_bottom_in[150], chany_bottom_in[156], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_30_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_30_sram_inv[0:11]),
		.out(chanx_left_out[154]));

	mux_2level_tapbuf_size28 mux_left_track_317 (
		.in({chany_top_in[1], chany_top_in[6], chany_top_in[55], chany_top_in[108], chanx_right_in[158], chany_bottom_in[51], chany_bottom_in[104], chany_bottom_in[154], chany_bottom_in[157], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_, left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_9_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_19_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_27_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_29_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_2_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.sram(mux_2level_tapbuf_size28_31_sram[0:11]),
		.sram_inv(mux_2level_tapbuf_size28_31_sram_inv[0:11]),
		.out(chanx_left_out[158]));

	mux_2level_tapbuf_size28_mem mem_left_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size29_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_0_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_0_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_77 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_1_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_1_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_2_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_2_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_3_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_3_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_101 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_4_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_4_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_109 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_5_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_5_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_117 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_6_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_6_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_125 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_7_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_7_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_133 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_8_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_8_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_141 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_9_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_9_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_149 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_10_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_10_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_157 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_11_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_11_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_165 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_12_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_12_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_173 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_13_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_13_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_181 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_14_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_14_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_189 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_15_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_15_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_197 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_16_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_16_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_205 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_17_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_17_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_213 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_18_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_18_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_221 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_19_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_19_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_229 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_20_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_20_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_237 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_21_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_21_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_245 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_22_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_22_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_253 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_23_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_23_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_261 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_24_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_24_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_269 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_25_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_25_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_277 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_26_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_26_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_285 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_27_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_27_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_293 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_28_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_28_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_301 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_29_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_29_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_309 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size28_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_30_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_30_sram_inv[0:11]));

	mux_2level_tapbuf_size28_mem mem_left_track_317 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size28_mem_30_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size28_31_sram[0:11]),
		.mem_outb(mux_2level_tapbuf_size28_31_sram_inv[0:11]));

endmodule
// ----- END Verilog module for sb_2__4_ -----

//----- Default net type -----
`default_nettype wire



