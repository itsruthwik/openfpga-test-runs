//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug 20 23:39:57 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__0_ -----
module sb_0__0_(pReset,
                prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:102] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:102] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:102] chany_top_out;
//----- OUTPUT PORTS -----
output [0:102] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_100_sram;
wire [0:1] mux_2level_tapbuf_size2_100_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_101_sram;
wire [0:1] mux_2level_tapbuf_size2_101_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_102_sram;
wire [0:1] mux_2level_tapbuf_size2_102_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_103_sram;
wire [0:1] mux_2level_tapbuf_size2_103_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_104_sram;
wire [0:1] mux_2level_tapbuf_size2_104_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_105_sram;
wire [0:1] mux_2level_tapbuf_size2_105_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_106_sram;
wire [0:1] mux_2level_tapbuf_size2_106_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_107_sram;
wire [0:1] mux_2level_tapbuf_size2_107_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_108_sram;
wire [0:1] mux_2level_tapbuf_size2_108_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_109_sram;
wire [0:1] mux_2level_tapbuf_size2_109_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_110_sram;
wire [0:1] mux_2level_tapbuf_size2_110_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_111_sram;
wire [0:1] mux_2level_tapbuf_size2_111_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_112_sram;
wire [0:1] mux_2level_tapbuf_size2_112_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_113_sram;
wire [0:1] mux_2level_tapbuf_size2_113_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_114_sram;
wire [0:1] mux_2level_tapbuf_size2_114_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_115_sram;
wire [0:1] mux_2level_tapbuf_size2_115_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_116_sram;
wire [0:1] mux_2level_tapbuf_size2_116_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_117_sram;
wire [0:1] mux_2level_tapbuf_size2_117_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_118_sram;
wire [0:1] mux_2level_tapbuf_size2_118_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_119_sram;
wire [0:1] mux_2level_tapbuf_size2_119_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_120_sram;
wire [0:1] mux_2level_tapbuf_size2_120_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_121_sram;
wire [0:1] mux_2level_tapbuf_size2_121_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_122_sram;
wire [0:1] mux_2level_tapbuf_size2_122_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_123_sram;
wire [0:1] mux_2level_tapbuf_size2_123_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_124_sram;
wire [0:1] mux_2level_tapbuf_size2_124_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_125_sram;
wire [0:1] mux_2level_tapbuf_size2_125_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_126_sram;
wire [0:1] mux_2level_tapbuf_size2_126_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_127_sram;
wire [0:1] mux_2level_tapbuf_size2_127_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_128_sram;
wire [0:1] mux_2level_tapbuf_size2_128_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_129_sram;
wire [0:1] mux_2level_tapbuf_size2_129_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_130_sram;
wire [0:1] mux_2level_tapbuf_size2_130_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_131_sram;
wire [0:1] mux_2level_tapbuf_size2_131_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_132_sram;
wire [0:1] mux_2level_tapbuf_size2_132_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_133_sram;
wire [0:1] mux_2level_tapbuf_size2_133_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_134_sram;
wire [0:1] mux_2level_tapbuf_size2_134_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_135_sram;
wire [0:1] mux_2level_tapbuf_size2_135_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_136_sram;
wire [0:1] mux_2level_tapbuf_size2_136_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_137_sram;
wire [0:1] mux_2level_tapbuf_size2_137_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_138_sram;
wire [0:1] mux_2level_tapbuf_size2_138_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_139_sram;
wire [0:1] mux_2level_tapbuf_size2_139_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_140_sram;
wire [0:1] mux_2level_tapbuf_size2_140_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_141_sram;
wire [0:1] mux_2level_tapbuf_size2_141_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_142_sram;
wire [0:1] mux_2level_tapbuf_size2_142_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_143_sram;
wire [0:1] mux_2level_tapbuf_size2_143_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_144_sram;
wire [0:1] mux_2level_tapbuf_size2_144_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_145_sram;
wire [0:1] mux_2level_tapbuf_size2_145_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_146_sram;
wire [0:1] mux_2level_tapbuf_size2_146_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_147_sram;
wire [0:1] mux_2level_tapbuf_size2_147_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_148_sram;
wire [0:1] mux_2level_tapbuf_size2_148_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_149_sram;
wire [0:1] mux_2level_tapbuf_size2_149_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_150_sram;
wire [0:1] mux_2level_tapbuf_size2_150_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_151_sram;
wire [0:1] mux_2level_tapbuf_size2_151_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_152_sram;
wire [0:1] mux_2level_tapbuf_size2_152_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_153_sram;
wire [0:1] mux_2level_tapbuf_size2_153_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_154_sram;
wire [0:1] mux_2level_tapbuf_size2_154_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_155_sram;
wire [0:1] mux_2level_tapbuf_size2_155_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_156_sram;
wire [0:1] mux_2level_tapbuf_size2_156_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_157_sram;
wire [0:1] mux_2level_tapbuf_size2_157_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_158_sram;
wire [0:1] mux_2level_tapbuf_size2_158_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_159_sram;
wire [0:1] mux_2level_tapbuf_size2_159_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_160_sram;
wire [0:1] mux_2level_tapbuf_size2_160_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_161_sram;
wire [0:1] mux_2level_tapbuf_size2_161_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_162_sram;
wire [0:1] mux_2level_tapbuf_size2_162_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_163_sram;
wire [0:1] mux_2level_tapbuf_size2_163_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_164_sram;
wire [0:1] mux_2level_tapbuf_size2_164_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_165_sram;
wire [0:1] mux_2level_tapbuf_size2_165_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_166_sram;
wire [0:1] mux_2level_tapbuf_size2_166_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_167_sram;
wire [0:1] mux_2level_tapbuf_size2_167_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_168_sram;
wire [0:1] mux_2level_tapbuf_size2_168_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_169_sram;
wire [0:1] mux_2level_tapbuf_size2_169_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_170_sram;
wire [0:1] mux_2level_tapbuf_size2_170_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_171_sram;
wire [0:1] mux_2level_tapbuf_size2_171_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_172_sram;
wire [0:1] mux_2level_tapbuf_size2_172_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_173_sram;
wire [0:1] mux_2level_tapbuf_size2_173_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_174_sram;
wire [0:1] mux_2level_tapbuf_size2_174_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_175_sram;
wire [0:1] mux_2level_tapbuf_size2_175_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_60_sram;
wire [0:1] mux_2level_tapbuf_size2_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_61_sram;
wire [0:1] mux_2level_tapbuf_size2_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_62_sram;
wire [0:1] mux_2level_tapbuf_size2_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_63_sram;
wire [0:1] mux_2level_tapbuf_size2_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_64_sram;
wire [0:1] mux_2level_tapbuf_size2_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_65_sram;
wire [0:1] mux_2level_tapbuf_size2_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_66_sram;
wire [0:1] mux_2level_tapbuf_size2_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_67_sram;
wire [0:1] mux_2level_tapbuf_size2_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_68_sram;
wire [0:1] mux_2level_tapbuf_size2_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_69_sram;
wire [0:1] mux_2level_tapbuf_size2_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_70_sram;
wire [0:1] mux_2level_tapbuf_size2_70_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_71_sram;
wire [0:1] mux_2level_tapbuf_size2_71_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_72_sram;
wire [0:1] mux_2level_tapbuf_size2_72_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_73_sram;
wire [0:1] mux_2level_tapbuf_size2_73_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_74_sram;
wire [0:1] mux_2level_tapbuf_size2_74_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_75_sram;
wire [0:1] mux_2level_tapbuf_size2_75_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_76_sram;
wire [0:1] mux_2level_tapbuf_size2_76_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_77_sram;
wire [0:1] mux_2level_tapbuf_size2_77_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_78_sram;
wire [0:1] mux_2level_tapbuf_size2_78_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_79_sram;
wire [0:1] mux_2level_tapbuf_size2_79_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_80_sram;
wire [0:1] mux_2level_tapbuf_size2_80_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_81_sram;
wire [0:1] mux_2level_tapbuf_size2_81_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_82_sram;
wire [0:1] mux_2level_tapbuf_size2_82_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_83_sram;
wire [0:1] mux_2level_tapbuf_size2_83_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_84_sram;
wire [0:1] mux_2level_tapbuf_size2_84_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_85_sram;
wire [0:1] mux_2level_tapbuf_size2_85_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_86_sram;
wire [0:1] mux_2level_tapbuf_size2_86_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_87_sram;
wire [0:1] mux_2level_tapbuf_size2_87_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_88_sram;
wire [0:1] mux_2level_tapbuf_size2_88_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_89_sram;
wire [0:1] mux_2level_tapbuf_size2_89_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_90_sram;
wire [0:1] mux_2level_tapbuf_size2_90_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_91_sram;
wire [0:1] mux_2level_tapbuf_size2_91_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_92_sram;
wire [0:1] mux_2level_tapbuf_size2_92_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_93_sram;
wire [0:1] mux_2level_tapbuf_size2_93_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_94_sram;
wire [0:1] mux_2level_tapbuf_size2_94_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_95_sram;
wire [0:1] mux_2level_tapbuf_size2_95_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_96_sram;
wire [0:1] mux_2level_tapbuf_size2_96_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_97_sram;
wire [0:1] mux_2level_tapbuf_size2_97_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_98_sram;
wire [0:1] mux_2level_tapbuf_size2_98_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_99_sram;
wire [0:1] mux_2level_tapbuf_size2_99_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:0] mux_2level_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_136_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_137_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_138_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_139_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_140_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_141_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_142_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_143_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_144_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_145_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_146_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_147_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_148_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_149_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_150_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_151_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_152_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_153_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_154_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_155_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_156_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_157_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_158_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_159_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_160_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_161_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_162_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_163_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_164_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_165_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_166_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_167_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_168_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_169_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_170_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_171_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_172_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_173_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_174_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_2level_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:0] mux_2level_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_2level_tapbuf_size3_mem_7_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chany_top_in[7];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chany_top_in[43];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[80] = chany_top_in[79];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chanx_right_in[9];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chanx_right_in[18];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chanx_right_in[27];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chanx_right_in[36];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chanx_right_in[45];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chanx_right_in[54];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chanx_right_in[63];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chanx_right_in[72];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chanx_right_in[81];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chanx_right_in[90];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chanx_right_in[99];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size3 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[1]}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_2level_tapbuf_size3 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[2]}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_2level_tapbuf_size3 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[3]}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_2level_tapbuf_size3 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[4]}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_2level_tapbuf_size3 mux_right_track_0 (
		.in({chany_top_in[102], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[0], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size3_mem mem_top_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_top_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[5]}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_2level_tapbuf_size2 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[6]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_2level_tapbuf_size2 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[7]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_2level_tapbuf_size2 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[8]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_2level_tapbuf_size2 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[10]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_2level_tapbuf_size2 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[11]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_2level_tapbuf_size2 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[12]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_2level_tapbuf_size2 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[13]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_2level_tapbuf_size2 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[14]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_2level_tapbuf_size2 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[15]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_2level_tapbuf_size2 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[16]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_2level_tapbuf_size2 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[17]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_2level_tapbuf_size2 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[19]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_2level_tapbuf_size2 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[20]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_2level_tapbuf_size2 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[21]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_2level_tapbuf_size2 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[22]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_2level_tapbuf_size2 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[23]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_2level_tapbuf_size2 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[24]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_2level_tapbuf_size2 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[25]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_2level_tapbuf_size2 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[26]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_2level_tapbuf_size2 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[28]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_2level_tapbuf_size2 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[29]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_2level_tapbuf_size2 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[30]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_2level_tapbuf_size2 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[31]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_2level_tapbuf_size2 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[32]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_2level_tapbuf_size2 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[33]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_2level_tapbuf_size2 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[34]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_2level_tapbuf_size2 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[35]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_2level_tapbuf_size2 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[37]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_2level_tapbuf_size2 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[38]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_2level_tapbuf_size2 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[39]}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_2level_tapbuf_size2 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[40]}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_2level_tapbuf_size2 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[41]}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_2level_tapbuf_size2 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[42]}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_2level_tapbuf_size2 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[43]}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_2level_tapbuf_size2 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[44]}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_2level_tapbuf_size2 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[46]}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_2level_tapbuf_size2 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[47]}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_2level_tapbuf_size2 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[48]}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_2level_tapbuf_size2 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[49]}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_2level_tapbuf_size2 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[50]}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_2level_tapbuf_size2 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[51]}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_2level_tapbuf_size2 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[52]}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_2level_tapbuf_size2 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[53]}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_2level_tapbuf_size2 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[55]}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_2level_tapbuf_size2 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[56]}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_2level_tapbuf_size2 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[57]}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_2level_tapbuf_size2 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[58]}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_2level_tapbuf_size2 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[59]}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_2level_tapbuf_size2 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[60]}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_2level_tapbuf_size2 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[61]}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_2level_tapbuf_size2 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[62]}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_2level_tapbuf_size2 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[64]}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_2level_tapbuf_size2 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[65]}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_2level_tapbuf_size2 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[66]}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_2level_tapbuf_size2 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[67]}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_2level_tapbuf_size2 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[68]}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_2level_tapbuf_size2 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[69]}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_2level_tapbuf_size2 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[70]}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_2level_tapbuf_size2 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[71]}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_2level_tapbuf_size2 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[73]}),
		.sram(mux_2level_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_60_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_2level_tapbuf_size2 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[74]}),
		.sram(mux_2level_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_61_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_2level_tapbuf_size2 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[75]}),
		.sram(mux_2level_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_62_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_2level_tapbuf_size2 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[76]}),
		.sram(mux_2level_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_63_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_2level_tapbuf_size2 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[77]}),
		.sram(mux_2level_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_64_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_2level_tapbuf_size2 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[78]}),
		.sram(mux_2level_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_65_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_2level_tapbuf_size2 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[79]}),
		.sram(mux_2level_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_66_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_2level_tapbuf_size2 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[80]}),
		.sram(mux_2level_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_67_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_2level_tapbuf_size2 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[82]}),
		.sram(mux_2level_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_68_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_2level_tapbuf_size2 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[83]}),
		.sram(mux_2level_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_69_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_2level_tapbuf_size2 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[84]}),
		.sram(mux_2level_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_70_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_2level_tapbuf_size2 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[85]}),
		.sram(mux_2level_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_71_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_2level_tapbuf_size2 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[86]}),
		.sram(mux_2level_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_72_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_2level_tapbuf_size2 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[87]}),
		.sram(mux_2level_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_73_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_2level_tapbuf_size2 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[88]}),
		.sram(mux_2level_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_74_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_2level_tapbuf_size2 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[89]}),
		.sram(mux_2level_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_75_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_2level_tapbuf_size2 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[91]}),
		.sram(mux_2level_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_76_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_2level_tapbuf_size2 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[92]}),
		.sram(mux_2level_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_77_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_2level_tapbuf_size2 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[93]}),
		.sram(mux_2level_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_78_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_2level_tapbuf_size2 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[94]}),
		.sram(mux_2level_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_79_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_2level_tapbuf_size2 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[95]}),
		.sram(mux_2level_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_80_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_2level_tapbuf_size2 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[96]}),
		.sram(mux_2level_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_81_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_2level_tapbuf_size2 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[97]}),
		.sram(mux_2level_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_82_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_2level_tapbuf_size2 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[98]}),
		.sram(mux_2level_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_83_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_2level_tapbuf_size2 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[100]}),
		.sram(mux_2level_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_84_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_2level_tapbuf_size2 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[101]}),
		.sram(mux_2level_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_85_sram_inv[0:1]),
		.out(chany_top_out[100]));

	mux_2level_tapbuf_size2 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[102]}),
		.sram(mux_2level_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_86_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_2level_tapbuf_size2 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[0]}),
		.sram(mux_2level_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_87_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_2level_tapbuf_size2 mux_right_track_8 (
		.in({chany_top_in[3], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_88_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size2 mux_right_track_10 (
		.in({chany_top_in[4], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_89_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size2 mux_right_track_12 (
		.in({chany_top_in[5], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_90_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size2 mux_right_track_14 (
		.in({chany_top_in[6], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_91_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size2 mux_right_track_18 (
		.in({chany_top_in[8], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_92_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size2 mux_right_track_20 (
		.in({chany_top_in[9], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_93_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size2 mux_right_track_22 (
		.in({chany_top_in[10], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_94_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size2 mux_right_track_24 (
		.in({chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_95_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size2 mux_right_track_26 (
		.in({chany_top_in[12], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_96_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size2 mux_right_track_28 (
		.in({chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_97_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size2 mux_right_track_30 (
		.in({chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_98_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size2 mux_right_track_32 (
		.in({chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_99_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size2 mux_right_track_36 (
		.in({chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_100_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size2 mux_right_track_38 (
		.in({chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_101_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size2 mux_right_track_40 (
		.in({chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_102_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size2 mux_right_track_42 (
		.in({chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_103_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size2 mux_right_track_44 (
		.in({chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_104_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size2 mux_right_track_46 (
		.in({chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_105_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size2 mux_right_track_48 (
		.in({chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_106_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size2 mux_right_track_50 (
		.in({chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_107_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size2 mux_right_track_54 (
		.in({chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_108_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size2 mux_right_track_56 (
		.in({chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_109_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size2 mux_right_track_58 (
		.in({chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_110_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size2 mux_right_track_60 (
		.in({chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_111_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size2 mux_right_track_62 (
		.in({chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_112_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size2 mux_right_track_64 (
		.in({chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_113_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size2 mux_right_track_66 (
		.in({chany_top_in[32], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_114_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size2 mux_right_track_68 (
		.in({chany_top_in[33], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_115_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size2 mux_right_track_72 (
		.in({chany_top_in[35], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_116_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size2 mux_right_track_74 (
		.in({chany_top_in[36], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_117_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size2 mux_right_track_76 (
		.in({chany_top_in[37], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_118_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size2 mux_right_track_78 (
		.in({chany_top_in[38], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_119_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size2 mux_right_track_80 (
		.in({chany_top_in[39], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_120_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size2 mux_right_track_82 (
		.in({chany_top_in[40], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_121_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size2 mux_right_track_84 (
		.in({chany_top_in[41], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_122_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size2 mux_right_track_86 (
		.in({chany_top_in[42], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_123_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size2 mux_right_track_90 (
		.in({chany_top_in[44], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_124_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size2 mux_right_track_92 (
		.in({chany_top_in[45], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_125_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size2 mux_right_track_94 (
		.in({chany_top_in[46], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_126_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size2 mux_right_track_96 (
		.in({chany_top_in[47], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_127_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size2 mux_right_track_98 (
		.in({chany_top_in[48], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_128_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size2 mux_right_track_100 (
		.in({chany_top_in[49], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_129_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_2level_tapbuf_size2 mux_right_track_102 (
		.in({chany_top_in[50], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_130_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_2level_tapbuf_size2 mux_right_track_104 (
		.in({chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_131_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_2level_tapbuf_size2 mux_right_track_108 (
		.in({chany_top_in[53], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_132_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_2level_tapbuf_size2 mux_right_track_110 (
		.in({chany_top_in[54], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_133_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_2level_tapbuf_size2 mux_right_track_112 (
		.in({chany_top_in[55], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_134_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_2level_tapbuf_size2 mux_right_track_114 (
		.in({chany_top_in[56], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_135_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_2level_tapbuf_size2 mux_right_track_116 (
		.in({chany_top_in[57], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_136_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_136_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_2level_tapbuf_size2 mux_right_track_118 (
		.in({chany_top_in[58], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_137_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_137_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_2level_tapbuf_size2 mux_right_track_120 (
		.in({chany_top_in[59], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_138_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_138_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_2level_tapbuf_size2 mux_right_track_122 (
		.in({chany_top_in[60], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_139_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_139_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_2level_tapbuf_size2 mux_right_track_126 (
		.in({chany_top_in[62], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_140_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_140_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_2level_tapbuf_size2 mux_right_track_128 (
		.in({chany_top_in[63], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_141_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_141_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_2level_tapbuf_size2 mux_right_track_130 (
		.in({chany_top_in[64], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_142_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_142_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_2level_tapbuf_size2 mux_right_track_132 (
		.in({chany_top_in[65], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_143_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_143_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_2level_tapbuf_size2 mux_right_track_134 (
		.in({chany_top_in[66], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_144_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_144_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_2level_tapbuf_size2 mux_right_track_136 (
		.in({chany_top_in[67], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_145_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_145_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_2level_tapbuf_size2 mux_right_track_138 (
		.in({chany_top_in[68], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_146_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_146_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_2level_tapbuf_size2 mux_right_track_140 (
		.in({chany_top_in[69], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_147_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_147_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_2level_tapbuf_size2 mux_right_track_144 (
		.in({chany_top_in[71], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_148_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_148_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_2level_tapbuf_size2 mux_right_track_146 (
		.in({chany_top_in[72], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_149_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_149_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_2level_tapbuf_size2 mux_right_track_148 (
		.in({chany_top_in[73], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_150_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_150_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_2level_tapbuf_size2 mux_right_track_150 (
		.in({chany_top_in[74], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_151_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_151_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_2level_tapbuf_size2 mux_right_track_152 (
		.in({chany_top_in[75], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_152_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_152_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_2level_tapbuf_size2 mux_right_track_154 (
		.in({chany_top_in[76], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_153_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_153_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_2level_tapbuf_size2 mux_right_track_156 (
		.in({chany_top_in[77], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_154_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_154_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_2level_tapbuf_size2 mux_right_track_158 (
		.in({chany_top_in[78], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_155_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_155_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_2level_tapbuf_size2 mux_right_track_162 (
		.in({chany_top_in[80], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_156_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_156_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_2level_tapbuf_size2 mux_right_track_164 (
		.in({chany_top_in[81], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_157_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_157_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_2level_tapbuf_size2 mux_right_track_166 (
		.in({chany_top_in[82], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_158_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_158_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_2level_tapbuf_size2 mux_right_track_168 (
		.in({chany_top_in[83], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_159_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_159_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_2level_tapbuf_size2 mux_right_track_170 (
		.in({chany_top_in[84], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_160_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_160_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_2level_tapbuf_size2 mux_right_track_172 (
		.in({chany_top_in[85], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_161_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_161_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_2level_tapbuf_size2 mux_right_track_174 (
		.in({chany_top_in[86], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_162_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_162_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_2level_tapbuf_size2 mux_right_track_176 (
		.in({chany_top_in[87], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_163_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_163_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_2level_tapbuf_size2 mux_right_track_180 (
		.in({chany_top_in[89], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_164_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_164_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_2level_tapbuf_size2 mux_right_track_182 (
		.in({chany_top_in[90], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_165_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_165_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_2level_tapbuf_size2 mux_right_track_184 (
		.in({chany_top_in[91], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_166_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_166_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_2level_tapbuf_size2 mux_right_track_186 (
		.in({chany_top_in[92], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_167_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_167_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_2level_tapbuf_size2 mux_right_track_188 (
		.in({chany_top_in[93], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_168_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_168_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_2level_tapbuf_size2 mux_right_track_190 (
		.in({chany_top_in[94], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_169_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_169_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_2level_tapbuf_size2 mux_right_track_192 (
		.in({chany_top_in[95], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_170_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_170_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_2level_tapbuf_size2 mux_right_track_194 (
		.in({chany_top_in[96], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_171_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_171_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_2level_tapbuf_size2 mux_right_track_198 (
		.in({chany_top_in[98], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_172_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_172_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_2level_tapbuf_size2 mux_right_track_200 (
		.in({chany_top_in[99], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_173_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_173_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_2level_tapbuf_size2 mux_right_track_202 (
		.in({chany_top_in[100], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_174_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_174_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_2level_tapbuf_size2 mux_right_track_204 (
		.in({chany_top_in[101], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_175_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_175_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_2level_tapbuf_size2_mem mem_top_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_60_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_61_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_62_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_63_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_64_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_65_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_66_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_67_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_68_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_69_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_70_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_71_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_72_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_73_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_74_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_75_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_76_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_77_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_78_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_79_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_80_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_81_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_82_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_83_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_84_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_85_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_86_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_top_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_87_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_88_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_89_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_90_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_91_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_92_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_93_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_94_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_95_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_96_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_97_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_98_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_99_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_100_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_101_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_102_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_103_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_104_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_105_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_106_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_107_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_108_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_109_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_110_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_111_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_112_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_113_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_114_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_115_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_116_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_117_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_118_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_119_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_120_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_121_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_122_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_123_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_124_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_125_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_126_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_127_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_128_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_100 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_129_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_102 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_130_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_104 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_131_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_108 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_132_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_110 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_133_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_112 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_134_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_114 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_135_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_116 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_136_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_136_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_118 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_136_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_137_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_137_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_120 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_137_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_138_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_138_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_122 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_138_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_139_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_139_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_126 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_139_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_140_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_140_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_128 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_140_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_141_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_141_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_130 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_141_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_142_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_142_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_132 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_142_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_143_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_143_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_134 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_143_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_144_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_144_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_136 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_144_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_145_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_145_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_138 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_145_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_146_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_146_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_140 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_146_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_147_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_147_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_144 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_147_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_148_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_148_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_146 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_148_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_149_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_149_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_148 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_149_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_150_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_150_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_150 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_150_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_151_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_151_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_152 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_151_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_152_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_152_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_154 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_152_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_153_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_153_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_156 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_153_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_154_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_154_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_158 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_154_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_155_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_155_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_162 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_155_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_156_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_156_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_164 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_156_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_157_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_157_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_166 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_157_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_158_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_158_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_168 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_158_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_159_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_159_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_170 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_159_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_160_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_160_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_172 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_160_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_161_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_161_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_174 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_161_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_162_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_162_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_176 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_162_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_163_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_163_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_180 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_163_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_164_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_164_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_182 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_164_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_165_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_165_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_184 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_165_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_166_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_166_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_186 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_166_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_167_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_167_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_188 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_167_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_168_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_168_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_190 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_168_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_169_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_169_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_192 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_169_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_170_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_170_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_194 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_170_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_171_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_171_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_198 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_171_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_172_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_172_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_200 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_172_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_173_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_173_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_202 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_173_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_174_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_174_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_204 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_174_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_175_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_175_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__0_ -----

//----- Default net type -----
`default_nettype wire



